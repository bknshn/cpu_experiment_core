module minrt (
  output logic [31:0] mem_inst [9999:0]
);
assign mem_inst [9365:0]= {32'hffffffff,32'h03e00008,32'h6c010000,32'h03e00008,32'hc7c00000,32'hafc10000,32'h00220825,32'h00021600,32'h68020000,32'h3c020000,32'h00220825,32'h00021400,32'h68020000,32'h3c020000,32'h00220825,32'h00021200,32'h68020000,32'h3c020000,32'h68010000,32'h3c010000,32'h03e00008,32'h00220825,32'h00021600,32'h68020000,32'h3c020000,32'h00220825,32'h00021400,32'h68020000,32'h3c020000,32'h00220825,32'h00021200,32'h68020000,32'h3c020000,32'h68010000,32'h3c010000,32'h03e00008,32'h46000007,32'h0800246b,32'h23bd0001,32'h2042ffff,32'he7a00000,32'h03e00008,32'h14400002,32'h37a10000,32'h34220000,32'h08002463,32'h23bd0001,32'h2063ffff,32'hafa20000,32'h03e00008,32'h14600002,32'h37a10000,32'h34230000,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc40005,32'h8fc30004,32'h8fc20003,32'h20050002,32'h20010000,32'h8fdf0007,32'h23defff8,32'h03400009,32'h23de0008,32'h8f7a0000,32'hafdf0007,32'h8fdb0001,32'h8fc10004,32'h20030000,32'h20020000,32'h8fdf0007,32'h23defff8,32'h0c0023bb,32'h23de0008,32'hafdf0007,32'h2021ffff,32'h8c210000,32'h20210000,32'h34210047,32'h3c010000,32'h8fdf0007,32'h23defff8,32'h0c001045,32'h23de0008,32'hafdf0007,32'h8fc10006,32'h8fdf0007,32'h23defff8,32'h0c0002de,32'h23de0008,32'hafdf0007,32'h3442008a,32'h3c020000,32'h8fdf0007,32'h23defff8,32'h0c00041e,32'h23de0008,32'hafdf0007,32'hafc10006,32'h34210040,32'h3c010000,32'h8fdf0006,32'h23defff9,32'h0c0022a0,32'h23de0007,32'hafdf0006,32'h8fdf0006,32'h23defff9,32'h0c001d7f,32'h23de0007,32'hafdf0006,32'h8fdf0006,32'h23defff9,32'h03400009,32'h23de0007,32'h8f7a0000,32'hafdf0006,32'hafc10005,32'h8fdb0002,32'h8fdf0005,32'h23defffa,32'h0c00206f,32'h23de0006,32'hafdf0005,32'hafc10004,32'h8fdf0004,32'h23defffb,32'h0c00206f,32'h23de0005,32'hafdf0004,32'hafc10003,32'h8fdf0003,32'h23defffc,32'h0c00206f,32'h23de0004,32'hafdf0003,32'hafc40002,32'hafc50001,32'hafc30000,32'he4200000,32'h20210000,32'h342100d8,32'h3c010000,32'h46010003,32'hc0210000,32'hc4400000,32'h34420000,32'h3c020000,32'hacc20000,32'h20c60001,32'h20020040,32'hace20000,32'h20c70000,32'h34c600d6,32'h3c060000,32'h20020040,32'hacc20000,32'h20c60001,32'hace10000,32'h20c70000,32'h34c600d4,32'h3c060000,32'h8f650001,32'h8f640002,32'h8f630003,32'h03e00008,32'h03e00008,32'h03e00008,32'h0800234a,32'h8fc20001,32'h8fc10000,32'h143a0004,32'h201a0002,32'h080022de,32'h8fc20001,32'h8fc10000,32'h143a0004,32'h201a0001,32'h8fdf0002,32'h23defffd,32'h0c0003b7,32'h23de0003,32'hafdf0002,32'h8fc10001,32'h03e00008,32'h143a0002,32'h201a0000,32'h8fdf0002,32'h23defffd,32'h0c000095,32'h23de0003,32'hafdf0002,32'hc4210000,32'h34210030,32'h3c010000,32'h8fdf0002,32'h23defffd,32'h0c0003de,32'h23de0003,32'hafdf0002,32'h8fc10001,32'h143a0023,32'h201a0002,32'h8fdf0002,32'h23defffd,32'h0c0003ba,32'h23de0003,32'hafdf0002,32'h20410000,32'hafc20001,32'hafc10000,32'h8c420000,32'h00411020,32'h13800030,32'h0341e02a,32'h201a0000,32'h34420048,32'h3c020000,32'h03e00008,32'hac410000,32'h20420000,32'h8fc20000,32'h20210001,32'h8fc10002,32'h8fdf000d,32'h23defff2,32'h0c0022b0,32'h23de000e,32'hafdf000d,32'h8fc20001,32'h8fc10002,32'hc7c2000b,32'hc7c10009,32'hc7c00005,32'h460100c1,32'hc4210000,32'h20210002,32'h8fc10006,32'h46010002,32'hc7c10007,32'h46000802,32'hc7c1000c,32'h8fdf000d,32'h23defff2,32'h0c0003cb,32'h23de000e,32'hafdf000d,32'h20410000,32'he7c2000c,32'he7c0000b,32'h8fc20003,32'hc4420000,32'h34420017,32'h3c020000,32'h46020001,32'hc4420000,32'h20220001,32'h8fc10006,32'h46010002,32'hc7c10007,32'h46000802,32'hc7c1000a,32'h8fdf000b,32'h23defff4,32'h0c0003c7,32'h23de000c,32'hafdf000b,32'h20410000,32'he7c2000a,32'he7c00009,32'h8fc20003,32'hc4420000,32'h34420017,32'h3c020000,32'h46020001,32'hc4420000,32'h20220000,32'h8fc10006,32'h46010002,32'hc7c10007,32'h46000802,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003c3,32'h23de000a,32'hafdf0009,32'he7c10008,32'he7c00007,32'h8fc10003,32'hc4210000,32'h34210017,32'h3c010000,32'h8fdf0007,32'h23defff8,32'h0c000338,32'h23de0008,32'hafdf0007,32'hafc10006,32'h3421008a,32'h3c010000,32'h20220000,32'h8fdf0006,32'h23defff9,32'h0c0003cf,32'h23de0007,32'hafdf0006,32'he7c00005,32'h8fc10003,32'h46000801,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0003de,32'h23de0006,32'hafdf0005,32'h20410000,32'he7c00004,32'hafc20003,32'hafc40002,32'hafc10001,32'hafc30000,32'hc4a00000,32'h34a50030,32'h3c050000,32'h8c840000,32'h20640000,32'h346301e3,32'h3c030000,32'h20210001,32'h00010880,32'h03e00008,32'hac410000,32'h20420000,32'h8fc20000,32'h20210003,32'h8fc10001,32'h8fdf0009,32'h23defff6,32'h0c0022b0,32'h23de000a,32'hafdf0009,32'h20620000,32'h20410000,32'hc7c20007,32'hc7c10006,32'hc7c00004,32'hc4830000,32'h20840002,32'h8fc40005,32'h20630003,32'h8fc30002,32'h20220002,32'h8fc10001,32'h8fdf0009,32'h23defff6,32'h0c0022b0,32'h23de000a,32'hafdf0009,32'h20820000,32'h20410000,32'hc7c30008,32'hc7c10006,32'hc7c00004,32'hc4c20000,32'h20a60001,32'h8fc50005,32'h20640002,32'h8fc30002,32'h20220001,32'h8fc10001,32'h8fdf0009,32'h23defff6,32'h0c0022b0,32'h23de000a,32'hafdf0009,32'h20810000,32'he7c30008,32'h8fc40001,32'hc7c20007,32'hc7c00004,32'hc4810000,32'h20640000,32'h8fc30005,32'h20220001,32'h8fc10002,32'h460000c6,32'h8fdf0008,32'h23defff7,32'h0c002471,32'h23de0009,32'hafdf0008,32'h46010006,32'he7c00007,32'hc4410000,32'h20220002,32'h8fc10005,32'h8fdf0007,32'h23defff8,32'h0c002471,32'h23de0008,32'hafdf0007,32'h46010006,32'he7c00006,32'hc4410000,32'h20220001,32'h8fc10005,32'h8fdf0006,32'h23defff9,32'h0c002471,32'h23de0007,32'hafdf0006,32'h46010006,32'hafc10005,32'he7c00004,32'hc4410000,32'h20220000,32'h3421008a,32'h3c010000,32'h46000801,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0003de,32'h23de0005,32'hafdf0004,32'h20410000,32'he7c00003,32'hafc10002,32'hafc40001,32'hafc30000,32'hc4a00000,32'h34a50030,32'h3c050000,32'h8c840000,32'h20640000,32'h346301e3,32'h3c030000,32'h00010880,32'h03e00008,32'hac410000,32'h00431020,32'h8fc30000,32'h3442012f,32'h3c020000,32'h20210000,32'hac220000,32'h8fc20001,32'hac220001,32'h8fc20006,32'he4200002,32'hc7c00002,32'h23bd0003,32'h23a10000,32'h8fdf0007,32'h23defff8,32'h0c001045,32'h23de0008,32'hafdf0007,32'h8fc10006,32'h8fdf0007,32'h23defff8,32'h0c0002cc,32'h23de0008,32'hafdf0007,32'hc7c20003,32'hc7c10004,32'hc7c00005,32'h8fdf0007,32'h23defff8,32'h0c00041e,32'h23de0008,32'hafdf0007,32'hafc10006,32'h8fdf0006,32'h23defff9,32'h0c002227,32'h23de0007,32'hafdf0006,32'he7c10005,32'he7c20004,32'he7c30003,32'he7c00002,32'hafc20001,32'hafc10000,32'h0800228c,32'h20010004,32'h8fdf0000,32'h23deffff,32'h0c002200,32'h23de0001,32'hafdf0000,32'h20030000,32'h20020000,32'h20010009,32'h8fdf0000,32'h23deffff,32'h0c002254,32'h23de0001,32'hafdf0000,32'h20010004,32'h03e00008,32'h0800228c,32'h2021ffff,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c00227a,32'h23de0002,32'hafdf0001,32'h20620000,32'h20410000,32'hafc10000,32'h20030077,32'h8c420000,32'h00411020,32'h1380000f,32'h0341e02a,32'h201a0000,32'h344200eb,32'h3c020000,32'h03e00008,32'h0800227a,32'h8fc10000,32'h2022ffff,32'h8fc10001,32'h8fdf0002,32'h23defffd,32'h0c001045,32'h23de0003,32'hafdf0002,32'h20610000,32'hafc20001,32'hafc10000,32'h8c630000,32'h00221820,32'h1380000f,32'h0342e02a,32'h201a0000,32'h03e00008,32'h08002254,32'h2021ffff,32'h8fc10000,32'h8fdf0003,32'h23defffc,32'h0c002242,32'h23de0004,32'hafdf0003,32'h20620000,32'h20030076,32'h8c210000,32'h00620820,32'hac810000,32'h00622020,32'h8fc30001,32'h8fc20000,32'h8fdf0003,32'h23defffc,32'h0c002461,32'h23de0004,32'hafdf0003,32'h8fc10002,32'h20220000,32'h8fdf0003,32'h23defffc,32'h0c002227,32'h23de0004,32'hafdf0003,32'hafc30002,32'hafc20001,32'hafc10000,32'h20030078,32'h13800021,32'h0341e02a,32'h201a0000,32'h344200eb,32'h3c020000,32'h03e00008,32'h08002242,32'h20610000,32'h2042ffff,32'hac810000,32'h00622020,32'h8fc30000,32'h8fc20001,32'h8fdf0002,32'h23defffd,32'h0c002227,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc10000,32'h1380000f,32'h0342e02a,32'h201a0000,32'h03e00008,32'h20410000,32'hac410000,32'h8fc10000,32'hac410001,32'h23bd0002,32'h23a20000,32'h8fdf0001,32'h23defffe,32'h0c002461,32'h23de0002,32'hafdf0001,32'hafc20000,32'h8c210000,32'h20210000,32'h34210047,32'h3c010000,32'h20220000,32'h8fdf0000,32'h23deffff,32'h0c002469,32'h23de0001,32'hafdf0000,32'hc4400000,32'h34420032,32'h3c020000,32'h20010003,32'h03e00008,32'h08002200,32'h8fc10003,32'h20230004,32'h8fc10000,32'h20220000,32'h8fdf0004,32'h23defffb,32'h0c0002c4,32'h23de0005,32'hafdf0004,32'h20610000,32'hafc10003,32'h8fc30001,32'h20020002,32'h2021ffff,32'h8fc10002,32'h8fdf0003,32'h23defffc,32'h0c0021b1,32'h23de0004,32'hafdf0003,32'h20810000,32'hafc10002,32'hafc20001,32'hafc30000,32'h20040004,32'h46010001,32'hc4810000,32'h34840001,32'h3c040000,32'h46010002,32'hc4810000,32'h34840024,32'h3c040000,32'hc0200000,32'h13800024,32'h0341e02a,32'h201a0000,32'h03e00008,32'h080021b1,32'h8fc30003,32'h8fc10004,32'hc7c00001,32'h20220000,32'h8fdf0005,32'h23defffa,32'h0c0002c4,32'h23de0006,32'hafdf0005,32'h20610000,32'hafc10004,32'h8fc30002,32'h20020001,32'h2021ffff,32'h8fc10000,32'h8fdf0004,32'h23defffb,32'h0c0020b3,32'h23de0005,32'hafdf0004,32'h20a20000,32'h20410000,32'h20830000,32'h8fc50002,32'hc7c30001,32'h20640002,32'h8fc30003,32'hc4610000,32'h34630032,32'h3c030000,32'hc4600000,32'h34630032,32'h3c030000,32'h20020000,32'h46010080,32'hc4410000,32'h34420004,32'h3c020000,32'h46010002,32'hc4410000,32'h34420024,32'h3c020000,32'hc0200000,32'h8fc10000,32'h8fdf0004,32'h23defffb,32'h0c0020b3,32'h23de0005,32'hafdf0004,32'h461f0046,32'h46010006,32'h460000c6,32'h460307c6,32'h20810000,32'hafc30003,32'hafc20002,32'he7c00001,32'hafc10000,32'hc4a30000,32'h34a50032,32'h3c050000,32'hc4a10000,32'h34a50032,32'h3c050000,32'h20040000,32'h46020881,32'hc4820000,32'h34840001,32'h3c040000,32'h46020842,32'hc4820000,32'h34840024,32'h3c040000,32'hc0210000,32'h1380004c,32'h0341e02a,32'h201a0000,32'h080020b3,32'h8fc30000,32'h8fc20001,32'h8fc10017,32'hc7c30014,32'hc7c20013,32'hc7c00016,32'h46000046,32'h8fdf0018,32'h23deffe7,32'h0c002097,32'h23de0019,32'hafdf0018,32'hafc10017,32'he7c00016,32'hc7c10014,32'h20210001,32'h8fc10015,32'h8fdf0016,32'h23deffe9,32'h0c002097,32'h23de0017,32'hafdf0016,32'h46020046,32'h46010006,32'hafc10015,32'he7c30014,32'hafc20001,32'hafc30000,32'he7c20013,32'h080002cc,32'h8fc10012,32'hc7c20008,32'hc7c10007,32'h8fdf0013,32'h23deffec,32'h0c002471,32'h23de0014,32'hafdf0013,32'hafc10012,32'hc7c00006,32'h8fdf0012,32'h23deffed,32'h0c00041e,32'h23de0013,32'hafdf0012,32'h8c210000,32'h00410820,32'h8fc20009,32'h20210051,32'h8fc10000,32'h8fdf0012,32'h23deffed,32'h0c0002cc,32'h23de0013,32'hafdf0012,32'h8fc10010,32'hc7c20008,32'hc7c00011,32'h46000046,32'h8fdf0012,32'h23deffed,32'h0c002471,32'h23de0013,32'hafdf0012,32'h46010006,32'he7c00011,32'hc7c10006,32'h8fdf0011,32'h23deffee,32'h0c002471,32'h23de0012,32'hafdf0011,32'hafc10010,32'hc7c00007,32'h8fdf0010,32'h23deffef,32'h0c00041e,32'h23de0011,32'hafdf0010,32'h20410000,32'h8c420000,32'h00621020,32'h8fc30009,32'h20220029,32'h8fc10000,32'h8fdf0010,32'h23deffef,32'h0c0002cc,32'h23de0011,32'hafdf0010,32'h8fc1000d,32'hc7c1000f,32'hc7c0000e,32'h46000086,32'h8fdf0010,32'h23deffef,32'h0c002471,32'h23de0011,32'hafdf0010,32'h46010006,32'he7c0000f,32'hc7c10006,32'h8fdf000f,32'h23defff0,32'h0c002471,32'h23de0010,32'hafdf000f,32'h46010006,32'he7c0000e,32'hc7c10008,32'h8fdf000e,32'h23defff1,32'h0c002471,32'h23de000f,32'hafdf000e,32'hafc1000d,32'hc7c00007,32'h8fdf000d,32'h23defff2,32'h0c00041e,32'h23de000e,32'hafdf000d,32'h20410000,32'h8c420000,32'h00621020,32'h8fc30009,32'h20220001,32'h8fc10000,32'h8fdf000d,32'h23defff2,32'h0c0002cc,32'h23de000e,32'hafdf000d,32'h8fc1000b,32'hc7c1000c,32'hc7c00006,32'h46000086,32'h8fdf000d,32'h23defff2,32'h0c002471,32'h23de000e,32'hafdf000d,32'h46010006,32'he7c0000c,32'hc7c10008,32'h8fdf000c,32'h23defff3,32'h0c002471,32'h23de000d,32'hafdf000c,32'hafc1000b,32'hc7c00007,32'h8fdf000b,32'h23defff4,32'h0c00041e,32'h23de000c,32'hafdf000b,32'h20410000,32'h8c420000,32'h00621020,32'h8fc30009,32'h20220050,32'h8fc10000,32'h8fdf000b,32'h23defff4,32'h0c0002cc,32'h23de000c,32'hafdf000b,32'h8fc1000a,32'hc7c10006,32'hc7c00007,32'h46000086,32'h8fdf000b,32'h23defff4,32'h0c002471,32'h23de000c,32'hafdf000b,32'hafc1000a,32'hc7c00008,32'h8fdf000a,32'h23defff5,32'h0c00041e,32'h23de000b,32'hafdf000a,32'h20410000,32'h8c420000,32'h00621020,32'h8fc30009,32'h20220028,32'h8fc10000,32'h8fdf000a,32'h23defff5,32'h0c0002cc,32'h23de000b,32'hafdf000a,32'hc7c20006,32'hc7c10008,32'hc7c00007,32'h8fdf000a,32'h23defff5,32'h0c00041e,32'h23de000b,32'hafdf000a,32'h20610000,32'hafc10009,32'he7c20008,32'he7c10007,32'he7c00006,32'h8c630000,32'h00221820,32'h8fc20000,32'h8c210000,32'h00410820,32'h8fc20002,32'h8fc10001,32'h46001803,32'hc4230000,32'h34210030,32'h3c010000,32'h46001083,32'hc7c20003,32'h46000843,32'hc7c10004,32'h46000004,32'h46010000,32'hc4210000,32'h34210030,32'h3c010000,32'h46000800,32'hc7c10005,32'h8fdf0006,32'h23defff9,32'h0c0000bb,32'h23de0007,32'hafdf0006,32'h46010006,32'he7c00005,32'hc7c10003,32'h8fdf0005,32'h23defffa,32'h0c0000bb,32'h23de0006,32'hafdf0005,32'he7c00004,32'he7c10003,32'hafc40002,32'hafc20001,32'hafc30000,32'h138000dc,32'h0341e02a,32'h201a0005,32'h348400eb,32'h3c040000,32'h03e00008,32'h46010002,32'hc7c10000,32'h8fdf0002,32'h23defffd,32'h0c002086,32'h23de0003,32'hafdf0002,32'h46010002,32'hc7c10001,32'h8fdf0002,32'h23defffd,32'h0c000223,32'h23de0003,32'hafdf0002,32'h46020006,32'he7c10001,32'he7c00000,32'h46001083,32'hc4220000,32'h34210030,32'h3c010000,32'h46000004,32'h46020000,32'hc4220000,32'h34210004,32'h3c010000,32'h46000002,32'h03e00008,32'h46000803,32'hc7c10001,32'h8fdf0002,32'h23defffd,32'h0c0000e6,32'h23de0003,32'hafdf0002,32'h46010006,32'he7c00001,32'hc7c10000,32'h8fdf0001,32'h23defffe,32'h0c00016d,32'h23de0002,32'hafdf0001,32'he7c00000,32'h0800205c,32'h2042fffe,32'h8c420000,32'h20420000,32'h8fc20000,32'h8fdf0002,32'h23defffd,32'h0c002461,32'h23de0003,32'hafdf0002,32'h8fc10001,32'h20220000,32'h8fdf0002,32'h23defffd,32'h0c00200a,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc10000,32'h8c420000,32'h20220000,32'h342100d4,32'h3c010000,32'h03e00008,32'h00010820,32'h0800205c,32'h20610000,32'h2042ffff,32'hac810000,32'h00622020,32'h8fc30000,32'h8fc20001,32'h8fdf0002,32'h23defffd,32'h0c00200a,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc10000,32'h1380000f,32'h0342e02a,32'h201a0000,32'h03e00008,32'h20410000,32'hac410000,32'h8fc10000,32'hac410001,32'h8fc10001,32'hac410002,32'h8fc10002,32'hac410003,32'h8fc10003,32'hac410004,32'h8fc10004,32'hac410005,32'h8fc10005,32'hac410006,32'h8fc10006,32'hac410007,32'h23bd0008,32'h23a20000,32'h8fdf0007,32'h23defff8,32'h0c001fc6,32'h23de0008,32'hafdf0007,32'hafc10006,32'h8fdf0006,32'h23defff9,32'h0c002461,32'h23de0007,32'hafdf0006,32'h20620000,32'h20410000,32'hafc10005,32'h20030000,32'h20020001,32'h8fdf0005,32'h23defffa,32'h0c001fc6,32'h23de0006,32'hafdf0005,32'hafc10004,32'h8fdf0004,32'h23defffb,32'h0c001fc6,32'h23de0005,32'hafdf0004,32'hafc10003,32'h8fdf0003,32'h23defffc,32'h0c002461,32'h23de0004,32'hafdf0003,32'h20620000,32'h20410000,32'hafc10002,32'h20030000,32'h20020005,32'h8fdf0002,32'h23defffd,32'h0c002461,32'h23de0003,32'hafdf0002,32'h20620000,32'h20410000,32'hafc10001,32'h20030000,32'h20020005,32'h8fdf0001,32'h23defffe,32'h0c001fc6,32'h23de0002,32'hafdf0001,32'hafc10000,32'h8fdf0000,32'h23deffff,32'h0c002469,32'h23de0001,32'hafdf0000,32'hc4400000,32'h34420032,32'h3c020000,32'h20010003,32'h03e00008,32'h00020820,32'hac610000,32'h20430004,32'h8fc20000,32'h8fdf0001,32'h23defffe,32'h0c002469,32'h23de0002,32'hafdf0001,32'hc4600000,32'h34630032,32'h3c030000,32'h20010003,32'hac610000,32'h20430003,32'h8fc20000,32'h8fdf0001,32'h23defffe,32'h0c002469,32'h23de0002,32'hafdf0001,32'hc4600000,32'h34630032,32'h3c030000,32'h20010003,32'hac610000,32'h20430002,32'h8fc20000,32'h8fdf0001,32'h23defffe,32'h0c002469,32'h23de0002,32'hafdf0001,32'hc4600000,32'h34630032,32'h3c030000,32'h20010003,32'hac610000,32'h20430001,32'h8fc20000,32'h8fdf0001,32'h23defffe,32'h0c002469,32'h23de0002,32'hafdf0001,32'h20410000,32'hafc10000,32'hc4600000,32'h34630032,32'h3c030000,32'h20020003,32'h8fdf0000,32'h23deffff,32'h0c002461,32'h23de0001,32'hafdf0000,32'h20010005,32'h20220000,32'h8fdf0000,32'h23deffff,32'h0c002469,32'h23de0001,32'hafdf0000,32'hc4400000,32'h34420032,32'h3c020000,32'h20010003,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc40004,32'h8fc30002,32'h8fc20003,32'h8fc10007,32'h20250000,32'h8fdf0008,32'h23defff7,32'h0c0002c4,32'h23de0009,32'hafdf0008,32'h20610000,32'hafc10007,32'h8fc30001,32'h20020002,32'h20210001,32'h8fc10005,32'h8fdf0007,32'h23defff8,32'h03400009,32'h23de0008,32'h8f7a0000,32'hafdf0007,32'h8fdb0006,32'h8fc50002,32'h8fc40003,32'h8fc30004,32'h8fc20005,32'h20010000,32'h8fdf0007,32'h23defff8,32'h03400009,32'h23de0008,32'h8f7a0000,32'hafdf0007,32'h20fb0000,32'h20810000,32'h21020000,32'h20a30000,32'h20280001,32'h08001fa7,32'h13800002,32'h0101e02a,32'hafc60006,32'hafc10005,32'hafc20004,32'hafc30003,32'hafc40002,32'hafc50001,32'hafdb0000,32'h2108ffff,32'h8d080000,32'h21080001,32'h03e00008,32'h13800002,32'h0121e02a,32'h8d290000,32'h21090001,32'h350800d4,32'h3c080000,32'h8f670001,32'h8f660002,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc50005,32'h8fc40004,32'h8fc30001,32'h8fc20006,32'h20210001,32'h8fc10007,32'h8fdf0009,32'h23defff6,32'h0c001de1,32'h23de000a,32'hafdf0009,32'h8fdf0009,32'h23defff6,32'h03400009,32'h23de000a,32'h8f7a0000,32'hafdf0009,32'h8fdb0002,32'h8fc50005,32'h8fc40004,32'h8fc30001,32'h8fc20006,32'h8fc10007,32'h20060000,32'h08001f78,32'h8fdf0009,32'h23defff6,32'h03400009,32'h23de000a,32'h8f7a0000,32'hafdf0009,32'h20610000,32'h20820000,32'h8fdb0003,32'h20040000,32'h8c630000,32'h00411820,32'h8fc20004,32'h8fc10007,32'h143a0010,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c001cbc,32'h23de000a,32'hafdf0009,32'h8fc30005,32'h8fc20006,32'h8fc10007,32'h8fdf0009,32'h23defff6,32'h0c0002de,32'h23de000a,32'hafdf0009,32'h8fc10008,32'h20220000,32'h8fdf0009,32'h23defff6,32'h0c000401,32'h23de000a,32'hafdf0009,32'h21010000,32'hafc90008,32'hafc10007,32'hafc20006,32'hafc50005,32'hafc40004,32'hafc70003,32'hafc60002,32'hafc30001,32'hafdb0000,32'h8d080000,32'h00814020,32'h03e00008,32'h13800002,32'h0101e02a,32'h352900d1,32'h3c090000,32'h8d080000,32'h21080000,32'h350800d4,32'h3c080000,32'h8f670001,32'h8f660002,32'h03400008,32'h8f7a0000,32'h461f0046,32'h46010006,32'h46000086,32'h460207c6,32'h2042ffff,32'h8c420000,32'h20420000,32'h344200d4,32'h3c020000,32'h46030000,32'hc4430000,32'h20820002,32'h46030002,32'hc4430000,32'h20420002,32'h46031080,32'hc4a30000,32'h20850001,32'h46020082,32'hc4a20000,32'h20450001,32'h46020840,32'hc4a20000,32'h20850000,32'h348400e5,32'h3c040000,32'h46010042,32'hc4810000,32'h20440000,32'h344200e2,32'h3c020000,32'h46010002,32'hc0410000,32'h00441022,32'h8c840000,32'h20840001,32'h348400d6,32'h3c040000,32'hc4800000,32'h20840000,32'h348400d8,32'h3c040000,32'h8f7b0001,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0003,32'h8fc2000d,32'h8fc1000a,32'hc7c20000,32'hc7c10001,32'hc7c00002,32'h20230000,32'h8fdf000e,32'h23defff1,32'h0c0002c4,32'h23de000f,32'hafdf000e,32'h20610000,32'hafc1000d,32'h8fc30005,32'h20020001,32'h2021ffff,32'h8fc10009,32'h8fdf000d,32'h23defff2,32'h03400009,32'h23de000e,32'h8f7a0000,32'hafdf000d,32'h20610000,32'h20820000,32'h8fdb0004,32'h20040000,32'h8c630000,32'h00411820,32'h8fc2000a,32'h8fc10009,32'h8fdf000d,32'h23defff2,32'h0c000417,32'h23de000e,32'hafdf000d,32'h20610000,32'h20820000,32'h8fc40005,32'h8c630000,32'h00411820,32'h8fc2000a,32'h8fc10009,32'h8fdf000d,32'h23defff2,32'h0c0002de,32'h23de000e,32'hafdf000d,32'h8fc20006,32'h8fdf000d,32'h23defff2,32'h0c000401,32'h23de000e,32'hafdf000d,32'h20610000,32'h8c630000,32'h00411820,32'h8fc2000a,32'h8fc10009,32'h8fdf000d,32'h23defff2,32'h03400009,32'h23de000e,32'h8f7a0000,32'hafdf000d,32'h20a20000,32'h20830000,32'h8fdb0008,32'h8fc50007,32'hc4a10000,32'h34a50032,32'h3c050000,32'h8c840000,32'h00622020,32'h8fc3000a,32'h8fc20009,32'hc4400000,32'h34420030,32'h3c020000,32'h20010000,32'h8fdf000d,32'h23defff2,32'h0c0002de,32'h23de000e,32'hafdf000d,32'h8fc2000b,32'h8fc1000c,32'h8fdf000d,32'h23defff2,32'h0c0002da,32'h23de000e,32'hafdf000d,32'h8fc10006,32'h8fdf000d,32'h23defff2,32'h0c0002eb,32'h23de000e,32'hafdf000d,32'h21610000,32'h21020000,32'hafc7000c,32'hafc6000b,32'hafc1000a,32'hafc20009,32'hafc40008,32'hafcb0007,32'hafca0006,32'hafc30005,32'hafc50004,32'hafdb0003,32'he7c00002,32'he7c10001,32'he7c20000,32'h20080000,32'he5030000,32'h21680002,32'h460218c0,32'h460418c2,32'hc5040000,32'h21080002,32'he5240000,32'h21690001,32'h46012100,32'h46041902,32'hc5240000,32'h21090001,32'he5240000,32'h21690000,32'h46002100,32'h46041902,32'hc5240000,32'h21090000,32'h460418c2,32'hc1240000,32'h00494822,32'h8d290000,32'h21890000,32'hc5230000,32'h21290000,32'h1380008f,32'h0342e02a,32'h201a0000,32'h358c00d6,32'h3c0c0000,32'h356b00e8,32'h3c0b0000,32'h354a00d1,32'h3c0a0000,32'h352900d8,32'h3c090000,32'h350800df,32'h3c080000,32'h34e700d9,32'h3c070000,32'h34c60087,32'h3c060000,32'h8f650001,32'h8f640002,32'h03e00008,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc10005,32'h20220001,32'h8fc10004,32'h8fdf0008,32'h23defff7,32'h0c0002de,32'h23de0009,32'hafdf0008,32'h20620000,32'h8fc30003,32'h8c210000,32'h00220820,32'h8fc20004,32'h8fdf0008,32'h23defff7,32'h0c000410,32'h23de0009,32'hafdf0008,32'h8fc10005,32'h8fdf0008,32'h23defff7,32'h03400009,32'h23de0009,32'h8f7a0000,32'hafdf0008,32'h20820000,32'h20410000,32'h20230000,32'h8fdb0001,32'h8c210000,32'h00230820,32'h8c840000,32'h00832020,32'h8fc40007,32'h8fc30004,32'h8c420000,32'h00621020,32'h8fc30002,32'h8fc20006,32'h8fdf0008,32'h23defff7,32'h0c000404,32'h23de0009,32'hafdf0008,32'h20410000,32'hafc10007,32'h8fc20005,32'h8fdf0007,32'h23defff8,32'h0c00041b,32'h23de0008,32'hafdf0007,32'h8fc10005,32'h8fdf0007,32'h23defff8,32'h0c0002da,32'h23de0008,32'hafdf0007,32'h20410000,32'hafc10006,32'h8fc20003,32'h8fdf0006,32'h23defff9,32'h0c000413,32'h23de0007,32'hafdf0006,32'h8fc10005,32'h08001e58,32'h143a0002,32'h201a0000,32'h8c210000,32'h00220820,32'h8fc20004,32'h8fdf0006,32'h23defff9,32'h0c00040a,32'h23de0007,32'hafdf0006,32'h8fc10005,32'h13800053,32'h0341e02a,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c001cd6,32'h23de0007,32'hafdf0006,32'hafc10005,32'hafc20004,32'hafc50003,32'hafc40002,32'hafc30001,32'hafdb0000,32'h13800062,32'h285c0004,32'h34a500ce,32'h3c050000,32'h348400eb,32'h3c040000,32'h8f630001,32'h08001dd5,32'hc4200000,32'h20210002,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c001dd5,32'h23de0002,32'hafdf0001,32'hc4400000,32'h20220001,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c001dd5,32'h23de0002,32'hafdf0001,32'hafc10000,32'hc4400000,32'h20220000,32'h342100d1,32'h3c010000,32'h08002493,32'h200100ff,32'h08001de0,32'h20010000,32'h08001dde,32'h00010820,32'h13800003,32'h0341e02a,32'h201a0000,32'h13800008,32'h283c00ff,32'he0010000,32'h08002493,32'h2001000a,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010035,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010035,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010032,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010020,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010038,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010032,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010031,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010020,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010038,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010032,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010031,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h2001000a,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010036,32'h8fdf0000,32'h23deffff,32'h0c002493,32'h23de0001,32'hafdf0000,32'h20010050,32'h03e00008,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0001,32'h8fc50005,32'h8fc40006,32'h8fc30007,32'h8fc20000,32'h8fc10008,32'h20260001,32'h8fc10004,32'h8fdf0009,32'h23defff6,32'h0c001c09,32'h23de000a,32'hafdf0009,32'h8fc40005,32'h8fc30006,32'h8fc20007,32'h8fc10008,32'h08001d73,32'h143a0002,32'h201a0000,32'h8c210000,32'h00250820,32'h8fc50004,32'h8fdf0009,32'h23defff6,32'h0c00040a,32'h23de000a,32'hafdf0009,32'h8fc10002,32'h03400008,32'h8f7a0000,32'h8fdb0003,32'h8fc20004,32'h8c210000,32'h00410820,32'h8fc20006,32'h8fc10008,32'h143a0009,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c001ce0,32'h23de000a,32'hafdf0009,32'h8fc50004,32'h8fc40005,32'h8fc30006,32'h8fc20007,32'h8fc10008,32'h13800034,32'h0341e02a,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c001cd6,32'h23de000a,32'hafdf0009,32'h21010000,32'h20c20000,32'hafc10008,32'hafc30007,32'hafc40006,32'hafc50005,32'hafc60004,32'hafc70003,32'hafc80002,32'hafdb0001,32'hafc20000,32'h13800048,32'h28dc0004,32'h8d080000,32'h00814020,32'h8f670001,32'h03e00008,32'h20010000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'h14220003,32'h8fc20005,32'h8fdf0006,32'h23defff9,32'h0c001cd6,32'h23de0007,32'hafdf0006,32'h20620000,32'h8fc30003,32'h8c210000,32'h00610820,32'h8fc30000,32'h20210001,32'h8fc10001,32'h14220013,32'h8fc20005,32'h8fdf0006,32'h23defff9,32'h0c001cd6,32'h23de0007,32'hafdf0006,32'h20610000,32'h20a20000,32'h8fc50003,32'h8c630000,32'h00831820,32'h8fc40000,32'h2023ffff,32'h8fc10001,32'h14220024,32'h8fc20005,32'h8fdf0006,32'h23defff9,32'h0c001cd6,32'h23de0007,32'hafdf0006,32'h20610000,32'h20820000,32'h8fc40003,32'h8c630000,32'h00611820,32'h8fc30002,32'h8fc10001,32'h14220034,32'h8fc20005,32'h8fdf0006,32'h23defff9,32'h0c001cd6,32'h23de0007,32'hafdf0006,32'h20610000,32'h20820000,32'hafc10005,32'h8fc40003,32'h8c630000,32'h00621820,32'h8fc30004,32'h8fc20001,32'h8fdf0005,32'h23defffa,32'h0c001cd6,32'h23de0006,32'hafdf0005,32'h20c10000,32'h20a20000,32'hafc20004,32'hafc50003,32'hafc40002,32'hafc10001,32'hafc30000,32'h8cc60000,32'h00613020,32'h03e00008,32'h8c210000,32'h00220820,32'h8fc20000,32'h8fdf0001,32'h23defffe,32'h0c000407,32'h23de0002,32'hafdf0001,32'hafc20000,32'h03e00008,32'h20010001,32'h03e00008,32'h20010000,32'h13800003,32'h283c0000,32'h03e00008,32'h20010000,32'h13800003,32'h0043e02a,32'h20230001,32'h8c420000,32'h20620000,32'h03e00008,32'h20010000,32'h13800003,32'h285c0000,32'h03e00008,32'h20010000,32'h13800003,32'h0085e02a,32'h20450001,32'h8c840000,32'h20640001,32'h346300d4,32'h3c030000,32'h03e00008,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc10003,32'h20220001,32'h8fc10002,32'h8fdf0004,32'h23defffb,32'h03400009,32'h23de0005,32'h8f7a0000,32'hafdf0004,32'h8fdb0001,32'h8fc10003,32'h08001cb4,32'h143a0002,32'h201a0000,32'h8c210000,32'h00220820,32'h8fc20002,32'h8fdf0004,32'h23defffb,32'h0c00040a,32'h23de0005,32'hafdf0004,32'h8fc10003,32'h1380001b,32'h0341e02a,32'h201a0000,32'h8c210000,32'h00220820,32'h8fc20002,32'h8fdf0004,32'h23defffb,32'h0c000407,32'h23de0005,32'hafdf0004,32'hafc10003,32'hafc20002,32'hafc30001,32'hafdb0000,32'h1380002b,32'h285c0004,32'h8f630001,32'h08000395,32'h8fc30009,32'h342100d1,32'h3c010000,32'h8c220000,32'h00220820,32'h8fc20000,32'h8fdf000a,32'h23defff5,32'h0c00040d,32'h23de000b,32'hafdf000a,32'h8c210000,32'h00410820,32'h8fc20003,32'h8fc10002,32'h8fdf000a,32'h23defff5,32'h0c00036f,32'h23de000b,32'hafdf000a,32'h20610000,32'h8fc30009,32'h8c420000,32'h00411020,32'h8fc20008,32'h8fc10000,32'h8fdf000a,32'h23defff5,32'h0c00036f,32'h23de000b,32'hafdf000a,32'h20610000,32'h8fc30009,32'h8c420000,32'h00411020,32'h8fc20007,32'h8fc10000,32'h8fdf000a,32'h23defff5,32'h0c00036f,32'h23de000b,32'hafdf000a,32'h20610000,32'h8fc30009,32'h8c420000,32'h00411020,32'h8fc20006,32'h8fc10000,32'h8fdf000a,32'h23defff5,32'h0c00036f,32'h23de000b,32'hafdf000a,32'h20610000,32'h8fc30009,32'h8c420000,32'h00411020,32'h8fc20005,32'h8fc10000,32'h8fdf000a,32'h23defff5,32'h0c0002de,32'h23de000b,32'hafdf000a,32'h20810000,32'h20620000,32'hafc40009,32'hafc10008,32'h348400ce,32'h3c040000,32'h8c630000,32'h00621820,32'h8fc30004,32'h8fc20000,32'h8fdf0008,32'h23defff7,32'h0c000410,32'h23de0009,32'hafdf0008,32'h20610000,32'hafc10007,32'h8c630000,32'h00621820,32'h8fc30001,32'h8fc20002,32'h8fdf0007,32'h23defff8,32'h0c000410,32'h23de0008,32'hafdf0007,32'h20610000,32'hafc10006,32'h8c630000,32'h00831820,32'h8fc40003,32'h20430001,32'h8fc20002,32'h8fdf0006,32'h23defff9,32'h0c000410,32'h23de0007,32'hafdf0006,32'h20810000,32'hafc10005,32'h8c840000,32'h00622020,32'h8fc30003,32'h8fc20002,32'h8fdf0005,32'h23defffa,32'h0c000410,32'h23de0006,32'hafdf0005,32'h20610000,32'hafc10004,32'h8c630000,32'h00831820,32'h8fc40003,32'h2043ffff,32'h8fc20002,32'h8fdf0004,32'h23defffb,32'h0c000410,32'h23de0005,32'hafdf0004,32'h20410000,32'hafc30003,32'hafc10002,32'hafc40001,32'hafc50000,32'h8c420000,32'h00411020,32'h08000395,32'h8fc30006,32'h342100d1,32'h3c010000,32'h8c220000,32'h00410820,32'h8fc20007,32'h8fc10001,32'h8fdf0008,32'h23defff7,32'h03400009,32'h23de0009,32'h8f7a0000,32'hafdf0008,32'h20830000,32'h20620000,32'h8fdb0000,32'h8c840000,32'h00822020,32'h8fc40005,32'h8c630000,32'h00621820,32'h8fc30004,32'h8fc20001,32'h8fdf0008,32'h23defff7,32'h0c000413,32'h23de0009,32'hafdf0008,32'h8fc10002,32'h8fdf0008,32'h23defff7,32'h0c0002de,32'h23de0009,32'hafdf0008,32'h20810000,32'h20620000,32'hafc10007,32'hafc40006,32'h348400ce,32'h3c040000,32'h8c630000,32'h00621820,32'h8fc30003,32'h8fc20001,32'h8fdf0006,32'h23defff9,32'h0c00040d,32'h23de0007,32'hafdf0006,32'h20410000,32'hafc10005,32'h8fc20002,32'h8fdf0005,32'h23defffa,32'h0c000404,32'h23de0006,32'hafdf0005,32'h20410000,32'hafc10004,32'h8fc20002,32'h8fdf0004,32'h23defffb,32'h0c00041b,32'h23de0005,32'hafdf0004,32'h20410000,32'hafc10003,32'h8fc20002,32'h8fdf0003,32'h23defffc,32'h0c000410,32'h23de0004,32'hafdf0003,32'hafc10002,32'hafc20001,32'hafc30000,32'h8f630001,32'h03400008,32'h8f7a0000,32'h8fdb0002,32'h8fc30000,32'h8fc20001,32'h8c210000,32'h20210004,32'h8fc10003,32'h03e00008,32'h143a0002,32'h201a0004,32'h8fc10004,32'h8fdf0005,32'h23defffa,32'h03400009,32'h23de0006,32'h8f7a0000,32'hafdf0005,32'h20a30000,32'h20610000,32'h20820000,32'h8fdb0002,32'h8fc50000,32'h8fc40001,32'h8c630000,32'h20430003,32'h8fc20003,32'h08001baf,32'h143a0002,32'h201a0003,32'h8fc10004,32'h8fdf0005,32'h23defffa,32'h03400009,32'h23de0006,32'h8f7a0000,32'hafdf0005,32'h20a30000,32'h20610000,32'h20820000,32'h8fdb0002,32'h8fc50000,32'h8fc40001,32'h8c630000,32'h20430002,32'h8fc20003,32'h08001b9c,32'h143a0002,32'h201a0002,32'h8fc10004,32'h8fdf0005,32'h23defffa,32'h03400009,32'h23de0006,32'h8f7a0000,32'hafdf0005,32'h20a30000,32'h20610000,32'h20820000,32'h8fdb0002,32'h8fc50000,32'h8fc40001,32'h8c630000,32'h20430001,32'h8fc20003,32'h08001b89,32'h143a0002,32'h201a0001,32'h8fc10004,32'h8fdf0005,32'h23defffa,32'h03400009,32'h23de0006,32'h8f7a0000,32'hafdf0005,32'h20a10000,32'h8ca50000,32'h20850000,32'h08001b76,32'h143a0002,32'h201a0000,32'hafc10004,32'hafc40003,32'hafdb0002,32'hafc20001,32'hafc30000,32'h348400eb,32'h3c040000,32'h8f7b0001,32'h03400008,32'h8f7a0000,32'h8fdb0003,32'h8fc30000,32'h8fc20001,32'h8fc10002,32'h20040076,32'h8fdf0004,32'h23defffb,32'h0c0010cf,32'h23de0005,32'hafdf0004,32'h20610000,32'hafc40003,32'hafc10002,32'hafc20001,32'hafc30000,32'h8f640001,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0002,32'h8fc30000,32'h8fc20001,32'h8fc10005,32'h2024fffe,32'h8fc10004,32'h8fdf0007,32'h23defff8,32'h03400009,32'h23de0008,32'h8f7a0000,32'hafdf0007,32'h20410000,32'h8fdb0003,32'h46000803,32'hc7c10006,32'hc4800000,32'h34840003,32'h3c040000,32'h8c420000,32'h00621020,32'h8fc30005,32'h20220001,32'h8fc10004,32'h08001b47,32'h8fdf0007,32'h23defff8,32'h03400009,32'h23de0008,32'h8f7a0000,32'hafdf0007,32'h20610000,32'h8fdb0003,32'h46000803,32'hc7c10006,32'hc4800000,32'h34840002,32'h3c040000,32'h8c630000,32'h00411820,32'h8fc20005,32'h8fc10004,32'h143a0013,32'h201a0000,32'h8fdf0007,32'h23defff8,32'h0c0000a4,32'h23de0008,32'hafdf0007,32'he7c00006,32'h8fdf0006,32'h23defff9,32'h0c000338,32'h23de0007,32'hafdf0006,32'h8fc20001,32'h8fdf0006,32'h23defff9,32'h0c00041e,32'h23de0007,32'hafdf0006,32'h20c10000,32'hafc10005,32'hafc40004,32'hafc50003,32'hafdb0002,32'hafc20001,32'hafc30000,32'h8cc60000,32'h00243020,32'h13800049,32'h0344e02a,32'h201a0000,32'h8f650001,32'h03e00008,32'h08000356,32'h8fc20003,32'h8fc10004,32'h46000802,32'hc7c1000a,32'h8fdf000b,32'h23defff4,32'h0c0003de,32'h23de000c,32'hafdf000b,32'he7c0000a,32'h8fc10008,32'h46000802,32'hc7c10000,32'h46000006,32'hc7c00009,32'h08001af4,32'hc4200000,32'h34210032,32'h3c010000,32'h143a0005,32'h201a0000,32'h8fdf000a,32'h23defff5,32'h0c00009b,32'h23de000b,32'hafdf000a,32'he7c00009,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'h8fdf0009,32'h23defff6,32'h0c000338,32'h23de000a,32'hafdf0009,32'h8fc20005,32'h8fc10006,32'h143a0029,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c00126b,32'h23de000a,32'hafdf0009,32'h8c420000,32'h20420000,32'h8fc20001,32'h20010000,32'h8fdf0009,32'h23defff6,32'h0c001622,32'h23de000a,32'hafdf0009,32'h8fc20007,32'h8fc10008,32'h8fdf0009,32'h23defff6,32'h0c001611,32'h23de000a,32'hafdf0009,32'h8fc10008,32'h20220000,32'h8fdf0009,32'h23defff6,32'h0c00041e,32'h23de000a,32'hafdf0009,32'h20610000,32'hafc10008,32'hafc60007,32'hafc40006,32'hafc50005,32'hafc80004,32'hafc20003,32'h8fc30002,32'h8c210000,32'h00610820,32'h8c210000,32'h20e10000,32'h03e00008,32'h143a0002,32'h201a0000,32'h350800ce,32'h3c080000,32'h34e700c7,32'h3c070000,32'h34c600c4,32'h3c060000,32'h34a5008a,32'h3c050000,32'h348400c8,32'h3c040000,32'h34630048,32'h3c030000,32'h344200cb,32'h3c020000,32'h8fdf0003,32'h23defffc,32'h03400009,32'h23de0004,32'h8f7a0000,32'hafdf0003,32'hafc10002,32'hafc20001,32'he7c00000,32'h8f7b0001,32'h8f620002,32'h03e00008,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc30008,32'h8fc20012,32'h46011040,32'hc7c20001,32'hc4410000,32'h20420000,32'h8fc20002,32'h20210001,32'h8fc10013,32'h46000802,32'hc7c10010,32'h46000801,32'hc7c10020,32'h8fdf0021,32'h23deffde,32'h0c0003de,32'h23de0022,32'hafdf0021,32'h20410000,32'he7c00020,32'h8fc20018,32'hc4400000,32'h34420030,32'h3c020000,32'h145a001c,32'h201a0002,32'h8fc20019,32'hac430000,32'h00821020,32'h8fc40015,32'h2003ffff,32'h20220001,32'h08001a74,32'h13800002,32'h0341e02a,32'h201a0004,32'h8fc10013,32'h03e00008,32'h143a0002,32'h201a0000,32'h8fdf0020,32'h23deffdf,32'h0c000095,32'h23de0021,32'hafdf0020,32'hc7c10010,32'hc4200000,32'h34210004,32'h3c010000,32'h8fdf0020,32'h23deffdf,32'h03400009,32'h23de0021,32'h8f7a0000,32'hafdf0020,32'h8fdb0003,32'h8fc20012,32'hc7c1001e,32'hc7c0001a,32'h2021ffff,32'h8c210000,32'h20210000,32'h8fc10004,32'h8fdf0020,32'h23deffdf,32'h0c0010cf,32'h23de0021,32'hafdf0020,32'h8fc1000a,32'h08001a4a,32'h8fdf0020,32'h23deffdf,32'h0c001821,32'h23de0021,32'hafdf0020,32'hc7c2001e,32'hc7c0001f,32'h46000046,32'h8fdf0020,32'h23deffdf,32'h0c002471,32'h23de0021,32'hafdf0020,32'h8fdf0020,32'h23deffdf,32'h0c000338,32'h23de0021,32'hafdf0020,32'he7c0001f,32'h8fc20011,32'h8fc10012,32'h46010002,32'hc7c1001a,32'h8fdf001f,32'h23deffe0,32'h0c002471,32'h23de0020,32'hafdf001f,32'h8fdf001f,32'h23deffe0,32'h0c000338,32'h23de0020,32'hafdf001f,32'h8fc20011,32'h8fc10006,32'h143a0025,32'h201a0000,32'h8fdf001f,32'h23deffe0,32'h0c00126b,32'h23de0020,32'hafdf001f,32'he7c0001e,32'h8c420000,32'h20420000,32'h8fc20005,32'h20010000,32'h46000802,32'hc7c10010,32'h8fdf001e,32'h23deffe1,32'h0c0003e2,32'h23de001f,32'hafdf001e,32'h8fc10018,32'h8fdf001e,32'h23deffe1,32'h0c000356,32'h23de001f,32'hafdf001e,32'h8fc20006,32'h8fc10012,32'h46000802,32'hc7c1001d,32'h8fdf001e,32'h23deffe1,32'h0c000338,32'h23de001f,32'hafdf001e,32'he7c0001d,32'h8fc20006,32'h8fc10012,32'hc4200000,32'h34210005,32'h3c010000,32'hac610000,32'h00621820,32'h8fc3001b,32'h8fc20013,32'h20010000,32'h080019fe,32'h8fdf001d,32'h23deffe2,32'h0c0002de,32'h23de001e,32'hafdf001d,32'h20620000,32'h8fc30006,32'h8c210000,32'h00220820,32'h8fc20013,32'h8fdf001d,32'h23deffe2,32'h0c00041b,32'h23de001e,32'hafdf001d,32'h8fc10008,32'h8fdf001d,32'h23deffe2,32'h0c000385,32'h23de001e,32'hafdf001d,32'h20410000,32'h46010002,32'hc7c1001a,32'hc4600000,32'h34630006,32'h3c030000,32'h8c420000,32'h00411020,32'h8fc2001c,32'h8fc10013,32'h8fdf001d,32'h23deffe2,32'h0c0002de,32'h23de001e,32'hafdf001d,32'h20610000,32'h20820000,32'hafc1001c,32'h8fc40007,32'h8c630000,32'h00221820,32'h8fc20013,32'h8fdf001c,32'h23deffe3,32'h0c00040d,32'h23de001d,32'hafdf001c,32'h8fc10008,32'hac610000,32'h00621820,32'h8fc3001b,32'h8fc20013,32'h20010001,32'h143a0038,32'h201a0000,32'h8fdf001c,32'h23deffe3,32'h0c000095,32'h23de001d,32'hafdf001c,32'hc4210000,32'h34210031,32'h3c010000,32'h8fdf001c,32'h23deffe3,32'h0c0003de,32'h23de001d,32'hafdf001c,32'h20410000,32'hafc1001b,32'h8fc20018,32'h8fdf001b,32'h23deffe4,32'h0c00040a,32'h23de001c,32'hafdf001b,32'h8fc10008,32'h8fdf001b,32'h23deffe4,32'h0c0002de,32'h23de001c,32'hafdf001b,32'h20620000,32'h8fc3000a,32'h8c210000,32'h00220820,32'h8fc20013,32'h8fdf001b,32'h23deffe4,32'h0c000404,32'h23de001c,32'hafdf001b,32'h8fc10008,32'hac810000,32'h00622020,32'h8fc30015,32'h8fc20013,32'h00220820,32'h8c420000,32'h20420000,32'h8fc20009,32'h00010880,32'h8fc10017,32'h8fdf001b,32'h23deffe4,32'h0c001622,32'h23de001c,32'hafdf001b,32'h8fc2000a,32'h8fc10018,32'h8fdf001b,32'h23deffe4,32'h0c0002de,32'h23de001c,32'hafdf001b,32'h8fc2000a,32'h8fc1000b,32'h8fdf001b,32'h23deffe4,32'h0c001611,32'h23de001c,32'hafdf001b,32'he7c0001a,32'h8fc20012,32'h8fc10018,32'h46010002,32'hc7c10010,32'h8fdf001a,32'h23deffe5,32'h0c0003de,32'h23de001b,32'hafdf001a,32'h20410000,32'hafc10019,32'h8fc20018,32'h8fdf0019,32'h23deffe6,32'h0c0003ba,32'h23de001a,32'hafdf0019,32'h20410000,32'hafc20018,32'hafc10017,32'h8c420000,32'h00411020,32'h8fc2000c,32'h8c210000,32'h20210000,32'h8fc1000d,32'h03e00008,32'he4200000,32'h20210002,32'h46000800,32'hc4410000,32'h20220002,32'he4410000,32'h20220001,32'h46000840,32'hc4410000,32'h20220001,32'he4410000,32'h20220000,32'h46000840,32'hc4410000,32'h20220000,32'h8fc1000e,32'h46010002,32'hc4210000,32'h20210000,32'h8fc1000f,32'h46010002,32'hc7c10010,32'h46010002,32'hc7c10016,32'h8fdf0017,32'h23deffe8,32'h0c0000bb,32'h23de0018,32'hafdf0017,32'hc7c00016,32'h03e00008,32'h143a0002,32'h201a0000,32'h8fdf0017,32'h23deffe8,32'h0c00009b,32'h23de0018,32'hafdf0017,32'he7c00016,32'h8fdf0016,32'h23deffe9,32'h0c002471,32'h23de0017,32'hafdf0016,32'h8fdf0016,32'h23deffe9,32'h0c000338,32'h23de0017,32'hafdf0016,32'h8fc20011,32'h8fc10012,32'h03e00008,32'h145a0002,32'h201a0000,32'hac610000,32'h00621820,32'h8fc30015,32'h8fc20013,32'h2001ffff,32'h143a003d,32'h201a0000,32'h8fdf0016,32'h23deffe9,32'h03400009,32'h23de0017,32'h8f7a0000,32'hafdf0016,32'h20410000,32'hafc10015,32'h8fdb0014,32'h8fc20012,32'h8fdf0015,32'h23deffea,32'h0c000407,32'h23de0016,32'hafdf0015,32'h20610000,32'hafc60014,32'hafc10013,32'hafc20012,32'hafce0011,32'he7c00010,32'hafd2000f,32'hafca000e,32'hafd1000d,32'hafcb000c,32'hafc9000b,32'hafd0000a,32'hafcf0009,32'hafc30008,32'hafc80007,32'hafcc0006,32'hafc50005,32'hafcd0004,32'hafc40003,32'hafc70002,32'he7c10001,32'hafdb0000,32'h13800195,32'h283c0004,32'h3652008d,32'h3c120000,32'h363100c7,32'h3c110000,32'h361000c4,32'h3c100000,32'h35ef00c2,32'h3c0f0000,32'h35ce008a,32'h3c0e0000,32'h35ad01e3,32'h3c0d0000,32'h358c00c8,32'h3c0c0000,32'h356b0048,32'h3c0b0000,32'h354a00d1,32'h3c0a0000,32'h352900d9,32'h3c090000,32'h350800cb,32'h3c080000,32'h34e700c3,32'h3c070000,32'h8f660001,32'h8f650002,32'h8f640003,32'h03e00008,32'h03400008,32'h8f7a0000,32'h8fdb0000,32'h8fc20003,32'hc7c10002,32'hc7c00004,32'h2021ffff,32'h8fc10001,32'h080018d9,32'h080018d8,32'h8fdf0010,32'h23deffef,32'h0c001821,32'h23de0011,32'hafdf0010,32'hc7c20002,32'hc7c0000e,32'h46000842,32'hc7c1000f,32'h8fdf0010,32'h23deffef,32'h0c000338,32'h23de0011,32'hafdf0010,32'h8fc10003,32'h20220000,32'h8fdf0010,32'h23deffef,32'h0c00041e,32'h23de0011,32'hafdf0010,32'he7c0000f,32'he7c2000e,32'h8fc1000b,32'h46031082,32'hc7c3000d,32'h46010082,32'hc7c10004,32'h8fdf000e,32'h23defff1,32'h0c00042a,32'h23de000f,32'hafdf000e,32'he7c0000d,32'h8fc10007,32'h8fdf000d,32'h23defff2,32'h0c000338,32'h23de000e,32'hafdf000d,32'h8fc10005,32'h20220000,32'h8fdf000d,32'h23defff2,32'h0c00041e,32'h23de000e,32'hafdf000d,32'h8fc1000b,32'h143a0032,32'h201a0000,32'h8fdf000d,32'h23defff2,32'h0c00126b,32'h23de000e,32'hafdf000d,32'h8c420000,32'h20420000,32'h8fc20006,32'h20010000,32'h1441003e,32'h8fc2000c,32'h8fdf000d,32'h23defff2,32'h0c000424,32'h23de000e,32'hafdf000d,32'h20410000,32'hafc1000c,32'h8fc20007,32'h00220820,32'h8c420000,32'h20420000,32'h8fc20008,32'h00010880,32'h8c210000,32'h20210000,32'h8fc10009,32'h080018d9,32'h143a0002,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h03400009,32'h23de000d,32'h8f7a0000,32'hafdf000c,32'hafc1000b,32'h8fdb000a,32'h8fdf000b,32'h23defff4,32'h0c000427,32'h23de000c,32'hafdf000b,32'h20a10000,32'hafc4000a,32'hafc80009,32'hafc70008,32'hafc50007,32'hafc30006,32'hafc60005,32'he7c00004,32'hafc20003,32'he7c10002,32'hafc10001,32'hafdb0000,32'h8ca50000,32'h00a12820,32'h13800076,32'h0341e02a,32'h201a0000,32'h350800c7,32'h3c080000,32'h34e700c2,32'h3c070000,32'h34c600c8,32'h3c060000,32'h34a5012f,32'h3c050000,32'h8f640001,32'h8f630002,32'h03e00008,32'he4200000,32'h20210002,32'h46000800,32'hc4410000,32'h20220002,32'he4410000,32'h20220001,32'h46000840,32'hc4410000,32'h20220001,32'he4410000,32'h20220000,32'h46000840,32'hc4410000,32'h20220000,32'h8fc10003,32'h46010002,32'hc7c10000,32'h8fdf0004,32'h23defffb,32'h0c0000bb,32'h23de0005,32'hafdf0004,32'h8fdf0004,32'h23defffb,32'h0c0000bb,32'h23de0005,32'hafdf0004,32'hc7c00001,32'h03e00008,32'h143a0002,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c00009b,32'h23de0005,32'hafdf0004,32'hc7c00001,32'h8fdf0004,32'h23defffb,32'h0c000356,32'h23de0005,32'hafdf0004,32'h20610000,32'hc7c00002,32'h08001838,32'h143a0002,32'h201a0000,32'hafc30003,32'h346300d1,32'h3c030000,32'h344200cb,32'h3c020000,32'h8fdf0003,32'h23defffc,32'h0c00009b,32'h23de0004,32'hafdf0003,32'he7c00002,32'he7c10001,32'he7c20000,32'h03e00008,32'h03e00008,32'he4200000,32'h20210002,32'h8fc10003,32'h46010003,32'hc4210000,32'h3421000b,32'h3c010000,32'h46000802,32'hc4210000,32'h3421000c,32'h3c010000,32'hc4200000,32'h34210032,32'h3c010000,32'h08001814,32'h46000006,32'hc7c00020,32'h143a0004,32'h201a0000,32'h8fdf0021,32'h23deffde,32'h0c0000a4,32'h23de0022,32'hafdf0021,32'he7c00020,32'h46000801,32'hc7c1001f,32'h8fdf0020,32'h23deffdf,32'h0c0000bb,32'h23de0021,32'hafdf0020,32'h46010006,32'he7c0001f,32'h46020841,32'hc7c2001d,32'hc4210000,32'h34210031,32'h3c010000,32'h46000801,32'hc7c1001e,32'h8fdf001f,32'h23deffe0,32'h0c0000bb,32'h23de0020,32'hafdf001f,32'h46020006,32'he7c1001e,32'he7c0001d,32'h46031081,32'hc7c30018,32'hc4220000,32'h34210031,32'h3c010000,32'hc4210000,32'h3421000d,32'h3c010000,32'h46000801,32'hc7c1001c,32'h8fdf001d,32'h23deffe2,32'h0c000292,32'h23de001e,32'hafdf001d,32'he7c0001c,32'hc4200000,32'h34210010,32'h3c010000,32'h080017de,32'h46010003,32'hc4210000,32'h3421000e,32'h3c010000,32'h46010002,32'hc4210000,32'h3421000f,32'h3c010000,32'h8fdf001c,32'h23deffe3,32'h0c000223,32'h23de001d,32'hafdf001c,32'h46000005,32'h46000803,32'hc7c1001b,32'hc7c00016,32'h143a0013,32'h201a0000,32'h8fdf001c,32'h23deffe3,32'h0c000095,32'h23de001d,32'hafdf001c,32'h46020006,32'h46030046,32'he7c0001b,32'hc4230000,32'h34210011,32'h3c010000,32'h46010085,32'hc7c10016,32'h46000802,32'hc7c1001a,32'h46000004,32'h8fdf001b,32'h23deffe4,32'h0c0003c7,32'h23de001c,32'hafdf001b,32'he7c0001a,32'h8fc10001,32'h46000801,32'hc7c10019,32'h8fdf001a,32'h23deffe5,32'h0c0003d6,32'h23de001b,32'hafdf001a,32'he7c10019,32'he7c00018,32'h8fc10001,32'hc4210000,32'h20210001,32'h8fc10000,32'h46000801,32'hc7c10017,32'h8fdf0018,32'h23deffe7,32'h0c000292,32'h23de0019,32'hafdf0018,32'he7c00017,32'hc4200000,32'h34210010,32'h3c010000,32'h0800179b,32'h46010003,32'hc4210000,32'h3421000e,32'h3c010000,32'h46010002,32'hc4210000,32'h3421000f,32'h3c010000,32'h8fdf0017,32'h23deffe8,32'h0c000223,32'h23de0018,32'hafdf0017,32'h46000005,32'h46000803,32'hc7c10014,32'hc7c00011,32'h143a0013,32'h201a0000,32'h8fdf0017,32'h23deffe8,32'h0c000095,32'h23de0018,32'hafdf0017,32'h46020006,32'h46030046,32'he7c00016,32'hc4230000,32'h34210011,32'h3c010000,32'h46010085,32'hc7c10011,32'h46000800,32'hc7c10015,32'h8fdf0016,32'h23deffe9,32'h0c0000bb,32'h23de0017,32'hafdf0016,32'h46010006,32'he7c00015,32'hc7c10014,32'h8fdf0015,32'h23deffea,32'h0c0000bb,32'h23de0016,32'hafdf0015,32'h46010006,32'he7c00014,32'hc7c10011,32'h46000802,32'hc7c10013,32'h46000004,32'h8fdf0014,32'h23deffeb,32'h0c0003cb,32'h23de0015,32'hafdf0014,32'he7c00013,32'h8fc10001,32'h46000801,32'hc7c10012,32'h8fdf0013,32'h23deffec,32'h0c0003da,32'h23de0014,32'hafdf0013,32'h20410000,32'he7c10012,32'he7c00011,32'h8fc20001,32'hc4410000,32'h20220002,32'h8fc10000,32'h46000802,32'hc7c10010,32'h46000004,32'h8fdf0011,32'h23deffee,32'h0c0003c3,32'h23de0012,32'hafdf0011,32'he7c00010,32'h8fc10001,32'h46000801,32'hc7c1000f,32'h8fdf0010,32'h23deffef,32'h0c0003d2,32'h23de0011,32'hafdf0010,32'h20610000,32'he7c0000f,32'h8fc30001,32'hc4600000,32'h20430000,32'h8fc20000,32'h145a00eb,32'h201a0004,32'h03e00008,32'he4200000,32'h20210002,32'h46010002,32'hc4410000,32'h3442000c,32'h3c020000,32'h46000801,32'hc4410000,32'h34420030,32'h3c020000,32'he4410000,32'h20220001,32'h8fc10003,32'h46010042,32'hc4210000,32'h3421000c,32'h3c010000,32'h8fdf000f,32'h23defff0,32'h0c0000bb,32'h23de0010,32'hafdf000f,32'h8fdf000f,32'h23defff0,32'h0c0000e6,32'h23de0010,32'hafdf000f,32'h46010002,32'hc4210000,32'h3421000e,32'h3c010000,32'h46000801,32'hc7c1000e,32'h8fdf000f,32'h23defff0,32'h0c000292,32'h23de0010,32'hafdf000f,32'he7c0000e,32'h46010003,32'hc4210000,32'h3421000a,32'h3c010000,32'h46000004,32'h46000800,32'hc7c1000d,32'h8fdf000e,32'h23defff1,32'h0c0000bb,32'h23de000f,32'hafdf000e,32'h46010006,32'he7c0000d,32'hc7c1000c,32'h8fdf000d,32'h23defff2,32'h0c0000bb,32'h23de000e,32'hafdf000d,32'h46010006,32'he7c0000c,32'hc7c1000a,32'h46000801,32'hc7c1000b,32'h8fdf000c,32'h23defff3,32'h0c0003da,32'h23de000d,32'hafdf000c,32'he7c1000b,32'he7c0000a,32'h8fc10001,32'hc4210000,32'h20210002,32'h8fc10000,32'h46000801,32'hc7c10009,32'h8fdf000a,32'h23defff5,32'h0c0003d2,32'h23de000b,32'hafdf000a,32'h20610000,32'he7c00009,32'h8fc30001,32'hc4600000,32'h20430000,32'h8fc20000,32'h145a005a,32'h201a0003,32'h03e00008,32'he4200000,32'h20210001,32'h46000802,32'h46001001,32'hc4420000,32'h34420030,32'h3c020000,32'hc4410000,32'h3442000c,32'h3c020000,32'he4410000,32'h20220000,32'h8fc10003,32'h46000842,32'hc4210000,32'h3421000c,32'h3c010000,32'h8fdf0009,32'h23defff6,32'h0c0000bb,32'h23de000a,32'hafdf0009,32'h8fdf0009,32'h23defff6,32'h0c00016d,32'h23de000a,32'hafdf0009,32'h46010002,32'hc4410000,32'h34420009,32'h3c020000,32'hc4400000,32'h20420001,32'h8fc20000,32'h145a0024,32'h201a0002,32'h03e00008,32'he4200000,32'h20210001,32'h8fc10003,32'hc4200000,32'h3421000c,32'h3c010000,32'h080016b0,32'hc4200000,32'h34210032,32'h3c010000,32'h143a0005,32'h201a0000,32'h080016b0,32'hc4200000,32'h34210032,32'h3c010000,32'h080016a6,32'hc4200000,32'h3421000c,32'h3c010000,32'h143a0005,32'h201a0000,32'h145a000b,32'h201a0000,32'h8fc20006,32'h8fdf0009,32'h23defff6,32'h0c000095,32'h23de000a,32'hafdf0009,32'hc4210000,32'h3421000a,32'h3c010000,32'h46000801,32'hc7c10008,32'h46010002,32'hc4210000,32'h34210007,32'h3c010000,32'h8fdf0009,32'h23defff6,32'h0c000292,32'h23de000a,32'hafdf0009,32'h46010006,32'he7c00008,32'h46010042,32'hc4210000,32'h34210008,32'h3c010000,32'h46000801,32'hc7c10007,32'h8fdf0008,32'h23defff7,32'h0c0003da,32'h23de0009,32'hafdf0008,32'h20410000,32'he7c00007,32'hafc10006,32'h8fc20001,32'hc4400000,32'h20420002,32'h8fc20000,32'h8fdf0006,32'h23defff9,32'h0c000095,32'h23de0007,32'hafdf0006,32'hc4210000,32'h3421000a,32'h3c010000,32'h46000801,32'hc7c10005,32'h46010002,32'hc4210000,32'h34210007,32'h3c010000,32'h8fdf0006,32'h23defff9,32'h0c000292,32'h23de0007,32'hafdf0006,32'h46010006,32'he7c00005,32'h46010042,32'hc4210000,32'h34210008,32'h3c010000,32'h46000801,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0003d2,32'h23de0006,32'hafdf0005,32'h20610000,32'he7c00004,32'h8fc30001,32'hc4600000,32'h20430000,32'h8fc20000,32'h145a0068,32'h201a0001,32'h8fc20002,32'he4400000,32'h20220002,32'h8fc10003,32'h8fdf0004,32'h23defffb,32'h0c0003ee,32'h23de0005,32'hafdf0004,32'h20410000,32'h8fc20001,32'he4400000,32'h20220001,32'h8fc10003,32'h8fdf0004,32'h23defffb,32'h0c0003ea,32'h23de0005,32'hafdf0004,32'h20410000,32'hafc10003,32'h8fc20001,32'he4400000,32'h20220000,32'h342100cb,32'h3c010000,32'h8fdf0003,32'h23defffc,32'h0c0003e6,32'h23de0004,32'hafdf0003,32'h20410000,32'hafc10002,32'h8fc20001,32'h8fdf0002,32'h23defffd,32'h0c0003b4,32'h23de0003,32'hafdf0002,32'hafc10001,32'hafc20000,32'h08001555,32'h8fc10000,32'h08001526,32'h8fc10000,32'h143a0003,32'h201a0002,32'h08001501,32'h8fc10001,32'h143a0003,32'h201a0001,32'h8fdf0002,32'h23defffd,32'h0c0003b7,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc10000,32'h080002eb,32'h8fc1000b,32'h20220000,32'h8fdf000f,32'h23defff0,32'h0c0003bd,32'h23de0010,32'hafdf000f,32'h8fc10000,32'he4400000,32'h20220002,32'h8fc1000b,32'h46000800,32'hc7c1000a,32'h8fdf000f,32'h23defff0,32'h0c0000b6,32'h23de0010,32'hafdf000f,32'h46000800,32'hc7c1000e,32'h46000802,32'hc7c10005,32'h8fdf000f,32'h23defff0,32'h0c0003f2,32'h23de0010,32'hafdf000f,32'he7c0000e,32'h8fc10000,32'h46000802,32'hc7c10003,32'h8fdf000e,32'h23defff1,32'h0c0003f6,32'h23de000f,32'hafdf000e,32'h20410000,32'h8fc20000,32'he4400000,32'h20220001,32'h8fc1000b,32'h46000800,32'hc7c10009,32'h8fdf000e,32'h23defff1,32'h0c0000b6,32'h23de000f,32'hafdf000e,32'h46000800,32'hc7c1000d,32'h46000802,32'hc7c10007,32'h8fdf000e,32'h23defff1,32'h0c0003f2,32'h23de000f,32'hafdf000e,32'he7c0000d,32'h8fc10000,32'h46000802,32'hc7c10003,32'h8fdf000d,32'h23defff2,32'h0c0003fa,32'h23de000e,32'hafdf000d,32'h20410000,32'h8fc20000,32'he4400000,32'h20220000,32'h8fc1000b,32'h46000800,32'hc7c10008,32'h8fdf000d,32'h23defff2,32'h0c0000b6,32'h23de000e,32'hafdf000d,32'h46001000,32'hc7c2000c,32'h46000802,32'hc7c10007,32'h8fdf000d,32'h23defff2,32'h0c0003f6,32'h23de000e,32'hafdf000d,32'he7c0000c,32'h8fc10000,32'h46000802,32'hc7c10005,32'h8fdf000c,32'h23defff3,32'h0c0003fa,32'h23de000d,32'hafdf000c,32'h8fc10000,32'h08001608,32'he4200000,32'hc7c0000a,32'h20410002,32'he4200000,32'hc7c00009,32'h20410001,32'he4200000,32'hc7c00008,32'h20410000,32'h143a000b,32'h201a0000,32'hafc2000b,32'h344200c8,32'h3c020000,32'h8fdf000b,32'h23defff4,32'h0c0003c0,32'h23de000c,32'hafdf000b,32'he7c0000a,32'h8fc10000,32'h46000802,32'hc7c10007,32'h8fdf000a,32'h23defff5,32'h0c0003cb,32'h23de000b,32'hafdf000a,32'he7c00009,32'h8fc10000,32'h46000802,32'hc7c10005,32'h8fdf0009,32'h23defff6,32'h0c0003c7,32'h23de000a,32'hafdf0009,32'he7c00008,32'h8fc10000,32'h46000802,32'hc7c10003,32'h8fdf0008,32'h23defff7,32'h0c0003c3,32'h23de0009,32'hafdf0008,32'he7c00007,32'h8fc10000,32'h46000801,32'hc7c10006,32'h8fdf0007,32'h23defff8,32'h0c0003da,32'h23de0008,32'hafdf0007,32'he7c10006,32'he7c00005,32'h8fc10000,32'hc4210000,32'h20210002,32'h8fc10001,32'h46000801,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0003d6,32'h23de0006,32'hafdf0005,32'h20410000,32'he7c10004,32'he7c00003,32'h8fc20000,32'hc4410000,32'h20220001,32'h8fc10001,32'h46000801,32'hc7c10002,32'h8fdf0003,32'h23defffc,32'h0c0003d2,32'h23de0004,32'hafdf0003,32'he7c00002,32'hafc20001,32'hafc10000,32'hc4600000,32'h20430000,32'h344200c4,32'h3c020000,32'h03e00008,32'he4200000,32'h20210002,32'h8fc10001,32'h8fdf0002,32'h23defffd,32'h0c002471,32'h23de0003,32'hafdf0002,32'h8fdf0002,32'h23defffd,32'h0c0003cb,32'h23de0003,32'hafdf0002,32'h20410000,32'h8fc20000,32'he4400000,32'h20220001,32'h8fc10001,32'h8fdf0002,32'h23defffd,32'h0c002471,32'h23de0003,32'hafdf0002,32'h8fdf0002,32'h23defffd,32'h0c0003c7,32'h23de0003,32'hafdf0002,32'h20410000,32'hafc10001,32'h8fc20000,32'he4400000,32'h20220000,32'h342100c8,32'h3c010000,32'h8fdf0001,32'h23defffe,32'h0c002471,32'h23de0002,32'hafdf0001,32'h8fdf0001,32'h23defffe,32'h0c0003c3,32'h23de0002,32'hafdf0001,32'hafc10000,32'h03e00008,32'he4200000,32'h00410820,32'h8fc20000,32'h8fc10003,32'h8fdf0004,32'h23defffb,32'h0c002471,32'h23de0005,32'hafdf0004,32'h8fdf0004,32'h23defffb,32'h0c0002a3,32'h23de0005,32'hafdf0004,32'hafc20003,32'hc4200000,32'h00610820,32'h8fc30001,32'h2021ffff,32'h2022ffff,32'h8fc10002,32'h8fdf0003,32'h23defffc,32'h0c0002da,32'h23de0004,32'hafdf0003,32'h20610000,32'hafc20002,32'hafc10001,32'hafc30000,32'h346300c8,32'h3c030000,32'h8c420000,32'h20420000,32'h344200c2,32'h3c020000,32'h08000095,32'hc7c00001,32'hc4210000,32'h34210012,32'h3c010000,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0002,32'h23defffd,32'h0c000095,32'h23de0003,32'hafdf0002,32'he7c10001,32'hc4200000,32'h34210014,32'h3c010000,32'hc4210000,32'h20210000,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c001498,32'h23de0002,32'hafdf0001,32'h20810000,32'h20230000,32'hafc30000,32'h8c420000,32'h20420000,32'h20040000,32'he4800000,32'h20640000,32'h346300c3,32'h3c030000,32'hc4600000,32'h34630013,32'h3c030000,32'h8f620001,32'h08001498,32'h8fc30000,32'h8fc20001,32'h20210001,32'h8fc10002,32'h8fdf0006,32'h23defff9,32'h0c00147f,32'h23de0007,32'hafdf0006,32'h8fc30000,32'h8fc20003,32'h20010001,32'h080014d4,32'h143a0002,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c000095,32'h23de0007,32'hafdf0006,32'hc4210000,32'h20210000,32'h8fc10004,32'hc4200000,32'h20210000,32'h8fc10005,32'h080014d4,32'h143a0002,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c000d67,32'h23de0007,32'hafdf0006,32'h20a10000,32'h20620000,32'hafc70005,32'hafc60004,32'hafc40003,32'h080014d4,32'h8fdf0003,32'h23defffc,32'h0c00147f,32'h23de0004,32'hafdf0003,32'h20a10000,32'h20820000,32'h20050001,32'h14ba000a,32'h201a0063,32'hafc10002,32'hafc20001,32'hafc30000,32'h03e00008,32'h14ba0002,32'h201affff,32'h34e700c1,32'h3c070000,32'h34c600c3,32'h3c060000,32'h8ca50000,32'h20850000,32'h8c840000,32'h00412020,32'h0800147f,32'h8fc30000,32'h8fc20001,32'h20210001,32'h8fc10002,32'h8fdf0003,32'h23defffc,32'h0c0013dd,32'h23de0004,32'hafdf0003,32'h20a10000,32'h20820000,32'hafc10002,32'hafc20001,32'hafc30000,32'h20050000,32'h8c840000,32'h00a42020,32'h03e00008,32'h149a0002,32'h201affff,32'h34a5008f,32'h3c050000,32'h8c840000,32'h00412020,32'h080013dd,32'h8fc30002,32'h8fc20000,32'h20210001,32'h8fc10001,32'hac220000,32'h8fc2000c,32'h20210000,32'h8fc10003,32'hac220000,32'h8fc2000a,32'h20210000,32'h8fc10004,32'h8fdf0012,32'h23deffed,32'h0c0002cc,32'h23de0013,32'hafdf0012,32'h8fc10005,32'hc7c2000e,32'hc7c1000f,32'hc7c00010,32'he4200000,32'hc7c00011,32'h20210000,32'h8fc10008,32'h0800147a,32'h143a0002,32'h201a0000,32'h8fdf0012,32'h23deffed,32'h0c0011bf,32'h23de0013,32'hafdf0012,32'h46030086,32'h46020046,32'h46010006,32'he7c00011,32'he7c10010,32'he7c2000f,32'he7c3000e,32'h8fc20000,32'h20010000,32'h460418c0,32'hc4240000,32'h20410002,32'h460018c2,32'hc4230000,32'h20210002,32'h46031080,32'hc4630000,32'h20430001,32'h46001082,32'hc4620000,32'h20230001,32'h46020840,32'hc4620000,32'h20430000,32'h8fc20006,32'h46000842,32'hc4410000,32'h20220000,32'h8fc10007,32'h46000800,32'hc7c1000d,32'hc4200000,32'h34210015,32'h3c010000,32'h0800147a,32'h143a0002,32'h201a0000,32'h8fdf000e,32'h23defff1,32'h0c000095,32'h23de000f,32'hafdf000e,32'hc7c0000d,32'hc4410000,32'h20220000,32'h8fc10008,32'h0800147a,32'h143a0002,32'h201a0000,32'h8fdf000e,32'h23defff1,32'h0c000095,32'h23de000f,32'hafdf000e,32'he7c1000d,32'hafc1000c,32'hc4400000,32'h34420032,32'h3c020000,32'hc4410000,32'h20420000,32'h8fc20009,32'h080013dd,32'h8fc30002,32'h8fc20000,32'h20210001,32'h8fc10001,32'h03e00008,32'h143a0002,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h0c0003bd,32'h23de000d,32'hafdf000c,32'h8c210000,32'h00410820,32'h8fc2000b,32'h8fc1000a,32'h143a0012,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h0c000d67,32'h23de000d,32'hafdf000c,32'h20810000,32'h21820000,32'hafc8000b,32'hafc4000a,32'hafc70009,32'hafc50008,32'hafc10007,32'hafc60006,32'hafca0005,32'hafcb0004,32'hafc90003,32'h8fcc0002,32'h03e00008,32'h149a0002,32'h201affff,32'h356b00c7,32'h3c0b0000,32'h354a00c4,32'h3c0a0000,32'h352900c2,32'h3c090000,32'h35080048,32'h3c080000,32'h34e700c1,32'h3c070000,32'h34c600dc,32'h3c060000,32'h34a500c3,32'h3c050000,32'h8c840000,32'h00622020,32'h8fc30000,32'h8fc20001,32'h8fdf0003,32'h23defffc,32'h0c00041e,32'h23de0004,32'hafdf0003,32'h20610000,32'hafc30002,32'hafc10001,32'hafc20000,32'h08000095,32'hc7c00001,32'hc4210000,32'h34210012,32'h3c010000,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0002,32'h23defffd,32'h0c000095,32'h23de0003,32'hafdf0002,32'he7c10001,32'hc4200000,32'h34210014,32'h3c010000,32'hc4210000,32'h20210000,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c001371,32'h23de0002,32'hafdf0001,32'h20810000,32'h20230000,32'hafc30000,32'h8c420000,32'h20420000,32'h20040000,32'he4800000,32'h20640000,32'h346300c3,32'h3c030000,32'hc4600000,32'h34630013,32'h3c030000,32'h8f620001,32'h08001371,32'h8fc30000,32'h8fc20001,32'h20210001,32'h8fc10002,32'h8fdf0006,32'h23defff9,32'h0c001358,32'h23de0007,32'hafdf0006,32'h8fc30000,32'h8fc20003,32'h20010001,32'h080013b0,32'h143a0002,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c000095,32'h23de0007,32'hafdf0006,32'hc4210000,32'h20210000,32'h8fc10004,32'hc4200000,32'h20210000,32'h8fc10005,32'h080013b0,32'h143a0002,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c000ab1,32'h23de0007,32'hafdf0006,32'h20e30000,32'h20a10000,32'h20620000,32'hafc80005,32'hafc60004,32'hafc40003,32'h080013b0,32'h8fdf0003,32'h23defffc,32'h0c001358,32'h23de0004,32'hafdf0003,32'h20a10000,32'h20820000,32'h20050001,32'h14ba000a,32'h201a0063,32'hafc10002,32'hafc20001,32'hafc30000,32'h03e00008,32'h14ba0002,32'h201affff,32'h350800c1,32'h3c080000,32'h34e700d9,32'h3c070000,32'h34c600c3,32'h3c060000,32'h8ca50000,32'h20850000,32'h8c840000,32'h00412020,32'h08001358,32'h8fc30000,32'h8fc20001,32'h20210001,32'h8fc10002,32'h8fdf0003,32'h23defffc,32'h0c0012bd,32'h23de0004,32'hafdf0003,32'h20a10000,32'h20820000,32'hafc10002,32'hafc20001,32'hafc30000,32'h20050000,32'h8c840000,32'h00a42020,32'h03e00008,32'h149a0002,32'h201affff,32'h34a5008f,32'h3c050000,32'h8c840000,32'h00412020,32'h080012bd,32'h8fc30006,32'h8fc20007,32'h20210001,32'h8fc10008,32'hac220000,32'h8fc2000b,32'h20210000,32'h8fc10000,32'hac220000,32'h8fc20009,32'h20210000,32'h8fc10001,32'h8fdf0011,32'h23deffee,32'h0c0002cc,32'h23de0012,32'hafdf0011,32'h8fc10002,32'hc7c2000d,32'hc7c1000e,32'hc7c0000f,32'he4200000,32'hc7c00010,32'h20210000,32'h8fc10004,32'h08001353,32'h143a0002,32'h201a0000,32'h8fdf0011,32'h23deffee,32'h0c0011bf,32'h23de0012,32'hafdf0011,32'h46030086,32'h46020046,32'h46010006,32'h20620000,32'h20410000,32'he7c00010,32'he7c1000f,32'he7c2000e,32'he7c3000d,32'h8fc30007,32'h20020000,32'h460418c0,32'hc4440000,32'h20420002,32'h460018c2,32'hc4630000,32'h20230002,32'h46031080,32'hc4630000,32'h20430001,32'h46001082,32'hc4620000,32'h20230001,32'h46020840,32'hc4620000,32'h20430000,32'h8fc20003,32'h46000842,32'hc4410000,32'h20220000,32'h8fc10006,32'h46000800,32'hc7c1000c,32'hc4200000,32'h34210015,32'h3c010000,32'h08001353,32'h143a0002,32'h201a0000,32'h8fdf000d,32'h23defff2,32'h0c000095,32'h23de000e,32'hafdf000d,32'hc7c0000c,32'hc4410000,32'h20220000,32'h8fc10004,32'h08001353,32'h143a0002,32'h201a0000,32'h8fdf000d,32'h23defff2,32'h0c000095,32'h23de000e,32'hafdf000d,32'he7c1000c,32'hafc1000b,32'hc4400000,32'h34420032,32'h3c020000,32'hc4410000,32'h20420000,32'h8fc20005,32'h080012bd,32'h8fc30006,32'h8fc20007,32'h20210001,32'h8fc10008,32'h03e00008,32'h143a0002,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c0003bd,32'h23de000c,32'hafdf000b,32'h8c210000,32'h00410820,32'h8fc2000a,32'h8fc10009,32'h143a0012,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c000ab1,32'h23de000c,32'hafdf000b,32'h20c30000,32'h20810000,32'h20620000,32'hafc8000a,32'hafc40009,32'hafc10008,32'hafc20007,32'hafc30006,32'hafc70005,32'hafc50004,32'hafc60003,32'hafca0002,32'hafcb0001,32'hafc90000,32'h03e00008,32'h149a0002,32'h201affff,32'h356b00c7,32'h3c0b0000,32'h354a00c4,32'h3c0a0000,32'h352900c2,32'h3c090000,32'h35080048,32'h3c080000,32'h34e700c1,32'h3c070000,32'h34c600d9,32'h3c060000,32'h34a500c3,32'h3c050000,32'h8c840000,32'h00412020,32'h03e00008,32'h20010001,32'h0800126b,32'h8fc20001,32'h20210001,32'h8fc10002,32'h143a0005,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c00124f,32'h23de0005,32'hafdf0004,32'h8fc20000,32'h20010001,32'h0800126b,32'h8fc20001,32'h20210001,32'h8fc10002,32'h143a0005,32'h201a0000,32'h20010001,32'h080012a8,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c00124f,32'h23de0005,32'hafdf0004,32'h8fc20000,32'h20010001,32'h080012a8,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c000095,32'h23de0005,32'hafdf0004,32'hc4210000,32'h34210014,32'h3c010000,32'hc4200000,32'h20210000,32'h8fc10003,32'h080012a8,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c000c92,32'h23de0005,32'hafdf0004,32'h20810000,32'h20c20000,32'h20e30000,32'hafc50003,32'h080012a8,32'h20010001,32'h149a0003,32'h201a0063,32'hafc10002,32'hafc20001,32'hafc30000,32'h03e00008,32'h20010000,32'h149a0003,32'h201affff,32'h34e700c4,32'h3c070000,32'h34c60040,32'h3c060000,32'h34a500c1,32'h3c050000,32'h8c840000,32'h20640000,32'h8c630000,32'h00411820,32'h03e00008,32'h20010001,32'h0800124f,32'h8fc20000,32'h20210001,32'h8fc10001,32'h143a0005,32'h201a0000,32'h8fdf0002,32'h23defffd,32'h0c0011df,32'h23de0003,32'hafdf0002,32'h20810000,32'h20620000,32'hafc10001,32'hafc20000,32'h20040000,32'h8c630000,32'h00831820,32'h03e00008,32'h20010000,32'h147a0003,32'h201affff,32'h3484008f,32'h3c040000,32'h8c630000,32'h00411820,32'h03e00008,32'h20010001,32'h080011df,32'h8fc20002,32'h20210001,32'h8fc10003,32'h143a0005,32'h201a0000,32'h8fdf0008,32'h23defff7,32'h0c0011bf,32'h23de0009,32'hafdf0008,32'h461f0046,32'h46010006,32'h46000086,32'h460207c6,32'h8fc20002,32'h20010000,32'h46030000,32'hc4230000,32'h20410002,32'h46001802,32'hc4230000,32'h20210002,32'h46031080,32'hc4630000,32'h20430001,32'h46001082,32'hc4620000,32'h20230001,32'h46020840,32'hc4620000,32'h20430000,32'h8fc20000,32'h46000842,32'hc4410000,32'h20220000,32'h8fc10001,32'h46000800,32'hc7c10007,32'hc4200000,32'h34210015,32'h3c010000,32'h080011df,32'h8fc20002,32'h20210001,32'h8fc10003,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0008,32'h23defff7,32'h0c0003bd,32'h23de0009,32'hafdf0008,32'h8c210000,32'h00410820,32'h8fc20005,32'h8fc10004,32'h143a0012,32'h201a0000,32'h8fdf0008,32'h23defff7,32'h0c000095,32'h23de0009,32'hafdf0008,32'hc4210000,32'h34210016,32'h3c010000,32'h08001210,32'h20010000,32'h143a0003,32'h201a0000,32'he7c00007,32'hc4400000,32'h20420000,32'h8fc20006,32'h8fdf0007,32'h23defff8,32'h0c000c92,32'h23de0008,32'hafdf0007,32'h21030000,32'h20610000,32'h20c20000,32'hafc40006,32'hafc50005,32'hafc30004,32'hafc10003,32'hafc20002,32'hafc70001,32'hafc80000,32'h8c630000,32'h00411820,32'h03e00008,32'h20010000,32'h147a0003,32'h201affff,32'h350800c4,32'h3c080000,32'h34e7008a,32'h3c070000,32'h34c60040,32'h3c060000,32'h34a50048,32'h3c050000,32'h348400c1,32'h3c040000,32'h8c630000,32'h00411820,32'h03e00008,32'h20010000,32'h080011bf,32'h8fc20003,32'hc7c20000,32'hc7c10001,32'hc7c00002,32'h20210001,32'h8fc10004,32'h143a0008,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c001188,32'h23de0006,32'hafdf0005,32'h20610000,32'hafc10004,32'hafc20003,32'he7c00002,32'he7c10001,32'he7c20000,32'h8c630000,32'h00831820,32'h03e00008,32'h20010001,32'h147a0003,32'h201affff,32'h34840048,32'h3c040000,32'h8c630000,32'h00411820,32'h08001156,32'h8fc10002,32'hc7c20006,32'hc7c10005,32'hc7c00004,32'h0800112a,32'h8fc10002,32'hc7c20006,32'hc7c10005,32'hc7c00004,32'h143a0006,32'h201a0002,32'h080010e1,32'h8fc10002,32'hc7c20006,32'hc7c10005,32'hc7c00004,32'h143a0006,32'h201a0001,32'h8fdf0007,32'h23defff8,32'h0c0003b7,32'h23de0008,32'hafdf0007,32'he7c00006,32'h8fc10002,32'h46000801,32'hc7c10000,32'h8fdf0006,32'h23defff9,32'h0c0003da,32'h23de0007,32'hafdf0006,32'he7c00005,32'h8fc10002,32'h46000801,32'hc7c10001,32'h8fdf0005,32'h23defffa,32'h0c0003d6,32'h23de0006,32'hafdf0005,32'he7c00004,32'h8fc10002,32'h46000801,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0003d2,32'h23de0005,32'hafdf0004,32'he7c00003,32'hafc10002,32'he7c10001,32'he7c20000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'h143a0003,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c000299,32'h23de0005,32'hafdf0004,32'h8fc10003,32'h20220000,32'h8fdf0004,32'h23defffb,32'h0c0000a4,32'h23de0005,32'hafdf0004,32'hafc10003,32'hc7c00002,32'h8fdf0003,32'h23defffc,32'h0c0003bd,32'h23de0004,32'hafdf0003,32'he7c00002,32'h8fc10000,32'h46000006,32'hc7c00001,32'h0800116d,32'h46000801,32'hc7c10001,32'hc4200000,32'h34210030,32'h3c010000,32'h143a0007,32'h201a0003,32'h8fdf0002,32'h23defffd,32'h0c0003b7,32'h23de0003,32'hafdf0002,32'he7c00001,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c000947,32'h23de0002,32'hafdf0001,32'hafc10000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'h143a0003,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c000299,32'h23de0007,32'hafdf0006,32'h8fc10005,32'h20220000,32'h8fdf0006,32'h23defff9,32'h0c0000a4,32'h23de0007,32'hafdf0006,32'hafc10005,32'hc7c00004,32'h8fdf0005,32'h23defffa,32'h0c0003bd,32'h23de0006,32'hafdf0005,32'he7c00004,32'h8fc10000,32'h8fdf0004,32'h23defffb,32'h0c00034a,32'h23de0005,32'hafdf0004,32'hc7c20001,32'hc7c10002,32'hc7c00003,32'h8fdf0004,32'h23defffb,32'h0c0003cf,32'h23de0005,32'hafdf0004,32'he7c00003,32'he7c10002,32'he7c20001,32'hafc10000,32'h080003bd,32'h8fc10001,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'h143a0003,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c0003bd,32'h23de0007,32'hafdf0006,32'h8fc10001,32'h143a000d,32'h201a0000,32'h8fdf0006,32'h23defff9,32'h0c000095,32'h23de0007,32'hafdf0006,32'hc7c00005,32'h46000046,32'h8fdf0006,32'h23defff9,32'h0c0003cb,32'h23de0007,32'hafdf0006,32'he7c00005,32'h8fc10001,32'h46000005,32'hc7c00000,32'h0800111a,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c000095,32'h23de0006,32'hafdf0005,32'hc7c00004,32'h46000046,32'h8fdf0005,32'h23defffa,32'h0c0003c7,32'h23de0006,32'hafdf0005,32'he7c00004,32'h8fc10001,32'h46000005,32'hc7c00002,32'h0800111a,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0004,32'h23defffb,32'h0c000095,32'h23de0005,32'hafdf0004,32'hc7c00003,32'h46000046,32'h8fdf0004,32'h23defffb,32'h0c0003c3,32'h23de0005,32'hafdf0004,32'he7c00003,32'he7c10002,32'hafc10001,32'he7c20000,32'h46000005,32'h0800104b,32'h8fc10000,32'h2022ffff,32'h8c210000,32'h20210000,32'h34210047,32'h3c010000,32'h8fdf0001,32'h23defffe,32'h0c0002de,32'h23de0002,32'hafdf0001,32'h23410000,32'h20220000,32'h205a0000,32'hafc10000,32'h344200dc,32'h3c020000,32'h03e00008,32'h0800104b,32'h8fc10002,32'h2022ffff,32'h8fc10000,32'he4200000,32'h20210003,32'h8fc10003,32'h46000006,32'h080010c7,32'h46010001,32'hc4210000,32'h34210030,32'h3c010000,32'h143a0006,32'h201a0003,32'h8fc10004,32'h8fdf0008,32'h23defff7,32'h0c000947,32'h23de0009,32'hafdf0008,32'h20610000,32'h8fc30001,32'hc4620000,32'h20230002,32'hc4610000,32'h20230001,32'hc4600000,32'h20230000,32'h080010ca,32'h13800002,32'h285c0002,32'h080010ca,32'he4200000,32'h20210003,32'h8fc10003,32'h8fdf0008,32'h23defff7,32'h0c00034a,32'h23de0009,32'hafdf0008,32'hc4620000,32'h20430002,32'hc4610000,32'h20430001,32'hc4600000,32'h20430000,32'h8fc20003,32'h8fdf0008,32'h23defff7,32'h0c0003cf,32'h23de0009,32'hafdf0008,32'h20410000,32'h8fc20001,32'h145a0018,32'h201a0002,32'h8fc20004,32'he4400000,32'h20220002,32'h8fc10003,32'h46000801,32'hc7c10007,32'h8fdf0008,32'h23defff7,32'h0c0003da,32'h23de0009,32'hafdf0008,32'h20610000,32'he7c00007,32'h8fc30001,32'hc4600000,32'h20430002,32'h8fc20002,32'he4400000,32'h20220001,32'h8fc10003,32'h46000801,32'hc7c10006,32'h8fdf0007,32'h23defff8,32'h0c0003d6,32'h23de0008,32'hafdf0007,32'h20610000,32'he7c00006,32'h8fc30001,32'hc4600000,32'h20430001,32'h8fc20002,32'he4400000,32'h20220000,32'h8fc10003,32'h46000801,32'hc7c10005,32'h8fdf0006,32'h23defff9,32'h0c0003d2,32'h23de0007,32'hafdf0006,32'h20610000,32'he7c00005,32'hafc10004,32'h8fc30001,32'hc4600000,32'h20430000,32'h8fc20002,32'h8fdf0004,32'h23defffb,32'h0c0003b7,32'h23de0005,32'hafdf0004,32'h20410000,32'hafc10003,32'h8fc20001,32'h8fdf0003,32'h23defffc,32'h0c0003fe,32'h23de0004,32'hafdf0003,32'h20610000,32'hafc10002,32'hafc30001,32'hafc20000,32'h8c630000,32'h00621820,32'h1380007f,32'h0342e02a,32'h201a0000,32'h34630048,32'h3c030000,32'h08000ffb,32'h2042ffff,32'h8c420000,32'h20420000,32'h34420047,32'h3c020000,32'h03e00008,32'h08000ffb,32'h8fc10000,32'h2042ffff,32'hac610000,32'h00621820,32'h8fc30003,32'h8fc20001,32'h8fdf0005,32'h23defffa,32'h0c000f06,32'h23de0006,32'hafdf0005,32'h8fc20002,32'h8fc10004,32'h08001041,32'hac610000,32'h00621820,32'h8fc30003,32'h8fc20001,32'h8fdf0005,32'h23defffa,32'h0c000e81,32'h23de0006,32'hafdf0005,32'h8fc20002,32'h8fc10004,32'h143a000d,32'h201a0002,32'h08001041,32'hac610000,32'h00621820,32'h8fc30003,32'h8fc20001,32'h8fdf0005,32'h23defffa,32'h0c000daf,32'h23de0006,32'hafdf0005,32'h8fc20002,32'h8fc10004,32'h143a000d,32'h201a0001,32'h8fdf0005,32'h23defffa,32'h0c0003b7,32'h23de0006,32'hafdf0005,32'h20410000,32'hafc10004,32'h8fc20002,32'h8fdf0004,32'h23defffb,32'h0c00041e,32'h23de0005,32'hafdf0004,32'h20410000,32'hafc10003,32'h8fc20000,32'h8fdf0003,32'h23defffc,32'h0c000421,32'h23de0004,32'hafdf0003,32'hafc30002,32'hafc20001,32'hafc10000,32'h8c630000,32'h00621820,32'h13800045,32'h0342e02a,32'h201a0000,32'h34630048,32'h3c030000,32'h03e00008,32'h00010820,32'h8fc10002,32'h08000ff8,32'he4400000,32'h20220004,32'h8fc10002,32'h46010003,32'hc7c10003,32'hc4200000,32'h34210030,32'h3c010000,32'h143a000a,32'h201a0000,32'h8fdf0013,32'h23deffec,32'h0c0000ad,32'h23de0014,32'hafdf0013,32'hc7c00003,32'he4400000,32'h20220003,32'h8fc10002,32'h46000801,32'hc7c10009,32'h8fdf0013,32'h23deffec,32'h0c0000b6,32'h23de0014,32'hafdf0013,32'h46000800,32'hc7c10011,32'h46000802,32'hc7c10012,32'h8fdf0013,32'h23deffec,32'h0c0003f6,32'h23de0014,32'hafdf0013,32'he7c10012,32'he7c00011,32'h8fc10000,32'hc4210000,32'h20210000,32'h8fc10001,32'h46000802,32'hc7c10010,32'h8fdf0011,32'h23deffee,32'h0c0003f2,32'h23de0012,32'hafdf0011,32'h20610000,32'he7c00010,32'h8fc30000,32'hc4600000,32'h20430001,32'h8fc20001,32'he4400000,32'h20220002,32'h8fc10002,32'h46000801,32'hc7c10007,32'h8fdf0010,32'h23deffef,32'h0c0000b6,32'h23de0011,32'hafdf0010,32'h46000800,32'hc7c1000e,32'h46000802,32'hc7c1000f,32'h8fdf0010,32'h23deffef,32'h0c0003fa,32'h23de0011,32'hafdf0010,32'h20410000,32'he7c1000f,32'he7c0000e,32'h8fc20000,32'hc4410000,32'h20220000,32'h8fc10001,32'h46000802,32'hc7c1000d,32'h8fdf000e,32'h23defff1,32'h0c0003f2,32'h23de000f,32'hafdf000e,32'h20610000,32'he7c0000d,32'h8fc30000,32'hc4600000,32'h20430002,32'h8fc20001,32'he4400000,32'h20220001,32'h8fc10002,32'h46000801,32'hc7c10005,32'h8fdf000d,32'h23defff2,32'h0c0000b6,32'h23de000e,32'hafdf000d,32'h46000800,32'hc7c1000b,32'h46000802,32'hc7c1000c,32'h8fdf000d,32'h23defff2,32'h0c0003fa,32'h23de000e,32'hafdf000d,32'h20410000,32'he7c1000c,32'he7c0000b,32'h8fc20000,32'hc4410000,32'h20220001,32'h8fc10001,32'h46000802,32'hc7c1000a,32'h8fdf000b,32'h23defff4,32'h0c0003f6,32'h23de000c,32'hafdf000b,32'h20410000,32'he7c0000a,32'h8fc20000,32'hc4400000,32'h20220002,32'h8fc10001,32'h08000fe7,32'he4400000,32'hc7c00009,32'h20220003,32'he4400000,32'hc7c00007,32'h20220002,32'he4400000,32'hc7c00005,32'h20220001,32'h8fc10002,32'h143a000c,32'h201a0000,32'h8fdf000a,32'h23defff5,32'h0c0003c0,32'h23de000b,32'hafdf000a,32'h20410000,32'he7c00009,32'h8fc20000,32'he4410000,32'hc7c10003,32'h20220000,32'h8fc10002,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'h46000802,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003cb,32'h23de000a,32'hafdf0009,32'h20410000,32'he7c10008,32'he7c00007,32'h8fc20000,32'hc4410000,32'h20220002,32'h8fc10001,32'h8fdf0007,32'h23defff8,32'h0c002471,32'h23de0008,32'hafdf0007,32'h46000802,32'hc7c10006,32'h8fdf0007,32'h23defff8,32'h0c0003c7,32'h23de0008,32'hafdf0007,32'h20410000,32'he7c10006,32'he7c00005,32'h8fc20000,32'hc4410000,32'h20220001,32'h8fc10001,32'h8fdf0005,32'h23defffa,32'h0c002471,32'h23de0006,32'hafdf0005,32'h46000802,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0003c3,32'h23de0006,32'hafdf0005,32'h20410000,32'he7c10004,32'he7c00003,32'h8fc20000,32'hc4410000,32'h20220000,32'h8fc10001,32'h8fdf0003,32'h23defffc,32'h0c000947,32'h23de0004,32'hafdf0003,32'h20610000,32'hafc10002,32'h8fc30000,32'hc4620000,32'h20430002,32'hc4610000,32'h20430001,32'hc4600000,32'h20430000,32'h8fc20001,32'h8fdf0002,32'h23defffd,32'h0c002469,32'h23de0003,32'hafdf0002,32'h20610000,32'hafc10001,32'hafc20000,32'hc4800000,32'h34840032,32'h3c040000,32'h20030005,32'h03e00008,32'h00010820,32'he4400000,32'h20220003,32'h8fc10002,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'h46010003,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003cb,32'h23de000a,32'hafdf0009,32'h20410000,32'h8fc20001,32'he4400000,32'h20220002,32'h8fc10002,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'h46010003,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003c7,32'h23de000a,32'hafdf0009,32'h20410000,32'h8fc20001,32'he4400000,32'h20220001,32'h8fc10002,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'h46010003,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003c3,32'h23de000a,32'hafdf0009,32'h20410000,32'h8fc20001,32'he4400000,32'h20220000,32'h8fc10002,32'h46010003,32'hc7c10008,32'hc4200000,32'h3421001b,32'h3c010000,32'h08000f04,32'he4400000,32'h20220000,32'h8fc10002,32'hc4200000,32'h34210032,32'h3c010000,32'h143a0008,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c00009b,32'h23de000a,32'hafdf0009,32'he7c00008,32'h46000800,32'hc7c10006,32'h46000802,32'hc7c10007,32'h8fdf0008,32'h23defff7,32'h0c0003cb,32'h23de0009,32'hafdf0008,32'he7c10007,32'he7c00006,32'h8fc10001,32'hc4210000,32'h20210002,32'h8fc10000,32'h46000800,32'hc7c10004,32'h46000802,32'hc7c10005,32'h8fdf0006,32'h23defff9,32'h0c0003c7,32'h23de0007,32'hafdf0006,32'h20410000,32'he7c10005,32'he7c00004,32'h8fc20001,32'hc4410000,32'h20220001,32'h8fc10000,32'h46000802,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0003c3,32'h23de0005,32'hafdf0004,32'h20610000,32'he7c00003,32'hafc10002,32'h8fc30001,32'hc4600000,32'h20430000,32'h8fc20000,32'h8fdf0002,32'h23defffd,32'h0c002469,32'h23de0003,32'hafdf0002,32'h20610000,32'hafc20001,32'hafc10000,32'hc4800000,32'h34840032,32'h3c040000,32'h20030004,32'h03e00008,32'h00010820,32'he4400000,32'h20220005,32'h8fc10002,32'hc4200000,32'h34210032,32'h3c010000,32'h08000e7f,32'he4400000,32'h20220005,32'h46010003,32'hc4410000,32'h20420002,32'h8fc20000,32'hc4400000,32'h34420030,32'h3c020000,32'he4400000,32'h20220004,32'h8fc10002,32'h8fdf0009,32'h23defff6,32'h0c0002bf,32'h23de000a,32'hafdf0009,32'h8fc10008,32'h8fdf0009,32'h23defff6,32'h0c0003cb,32'h23de000a,32'hafdf0009,32'h20410000,32'hafc10008,32'h8fc20001,32'h8fdf0008,32'h23defff7,32'h0c000299,32'h23de0009,32'hafdf0008,32'h8fc10007,32'h20220000,32'h8fdf0008,32'h23defff7,32'h0c0000a4,32'h23de0009,32'hafdf0008,32'hafc10007,32'hc4600000,32'h20430002,32'h8fc20000,32'h8fdf0007,32'h23defff8,32'h0c0003bd,32'h23de0008,32'hafdf0007,32'h8fc10001,32'h143a0032,32'h201a0000,32'h8fdf0007,32'h23defff8,32'h0c0000ad,32'h23de0008,32'hafdf0007,32'hc4600000,32'h20430002,32'h8fc20000,32'he4400000,32'h20220003,32'h8fc10002,32'hc4200000,32'h34210032,32'h3c010000,32'h08000e3e,32'he4600000,32'h20230003,32'h46010003,32'hc4610000,32'h20430001,32'h8fc20000,32'hc4400000,32'h34420030,32'h3c020000,32'he4400000,32'h20220002,32'h8fc10002,32'h8fdf0007,32'h23defff8,32'h0c0002bf,32'h23de0008,32'hafdf0007,32'h8fc10006,32'h8fdf0007,32'h23defff8,32'h0c0003c7,32'h23de0008,32'hafdf0007,32'h20410000,32'hafc10006,32'h8fc20001,32'h8fdf0006,32'h23defff9,32'h0c000299,32'h23de0007,32'hafdf0006,32'h8fc10005,32'h20220000,32'h8fdf0006,32'h23defff9,32'h0c0000a4,32'h23de0007,32'hafdf0006,32'hafc10005,32'hc4600000,32'h20430001,32'h8fc20000,32'h8fdf0005,32'h23defffa,32'h0c0003bd,32'h23de0006,32'hafdf0005,32'h8fc10001,32'h143a0032,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c0000ad,32'h23de0006,32'hafdf0005,32'hc4600000,32'h20430001,32'h8fc20000,32'he4400000,32'h20220001,32'h8fc10002,32'hc4200000,32'h34210032,32'h3c010000,32'h08000dfd,32'he4600000,32'h20230001,32'h46010003,32'hc4610000,32'h20430000,32'h8fc20000,32'hc4400000,32'h34420030,32'h3c020000,32'he4400000,32'h20220000,32'h8fc10002,32'h8fdf0005,32'h23defffa,32'h0c0002bf,32'h23de0006,32'hafdf0005,32'h8fc10004,32'h8fdf0005,32'h23defffa,32'h0c0003c3,32'h23de0006,32'hafdf0005,32'h20410000,32'hafc10004,32'h8fc20001,32'h8fdf0004,32'h23defffb,32'h0c000299,32'h23de0005,32'hafdf0004,32'h8fc10003,32'h20220000,32'h8fdf0004,32'h23defffb,32'h0c0000a4,32'h23de0005,32'hafdf0004,32'hafc10003,32'hc4600000,32'h20430000,32'h8fc20000,32'h8fdf0003,32'h23defffc,32'h0c0003bd,32'h23de0004,32'hafdf0003,32'h8fc10001,32'h143a0032,32'h201a0000,32'h8fdf0003,32'h23defffc,32'h0c0000ad,32'h23de0004,32'hafdf0003,32'hafc10002,32'hc4600000,32'h20430000,32'h8fc20000,32'h8fdf0002,32'h23defffd,32'h0c002469,32'h23de0003,32'hafdf0002,32'h20610000,32'hafc20001,32'hafc10000,32'hc4800000,32'h34840032,32'h3c040000,32'h20030006,32'h08000d09,32'h8fc30003,32'h8fc20007,32'h8fc10000,32'hc7c20004,32'hc7c10005,32'hc7c00006,32'h08000cef,32'h8fc30003,32'h8fc20007,32'h8fc10000,32'hc7c20004,32'hc7c10005,32'hc7c00006,32'h143a0008,32'h201a0002,32'h08000afa,32'h8fc30007,32'h8fc10000,32'hc7c20004,32'hc7c10005,32'hc7c00006,32'h20220000,32'h8fdf0008,32'h23defff7,32'h0c00041e,32'h23de0009,32'hafdf0008,32'h8fc10002,32'h143a000e,32'h201a0001,32'h8fdf0008,32'h23defff7,32'h0c0003b7,32'h23de0009,32'hafdf0008,32'h20410000,32'hafc10007,32'h8fc20000,32'h8c210000,32'h00220820,32'h8fc20001,32'h8fdf0007,32'h23defff8,32'h0c000421,32'h23de0008,32'hafdf0007,32'h20410000,32'he7c00006,32'he7c10005,32'he7c20004,32'hafc10003,32'h8fc20002,32'hc4420000,32'h20220002,32'hc4410000,32'h20220001,32'hc4400000,32'h20220000,32'h8fdf0003,32'h23defffc,32'h0c0003fe,32'h23de0004,32'hafdf0003,32'h20610000,32'hafc20002,32'hafc10001,32'hafc30000,32'h8c630000,32'h00611820,32'h34630048,32'h3c030000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'he4200000,32'h20210000,32'h8fc10007,32'h46010002,32'hc4210000,32'h20210004,32'h8fc10006,32'h46000800,32'hc7c10008,32'h46000004,32'hc7c0000a,32'h08000d63,32'he4200000,32'h20210000,32'h8fc10007,32'h46010002,32'hc4210000,32'h20210004,32'h8fc10006,32'h46000801,32'hc7c10008,32'h46000004,32'hc7c0000a,32'h143a000d,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c0003bd,32'h23de000c,32'hafdf000b,32'h8fc10000,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c00009b,32'h23de000c,32'hafdf000b,32'he7c0000a,32'h46010001,32'h46011042,32'hc7c20001,32'hc7c10009,32'h8fdf000a,32'h23defff5,32'h0c0000bb,32'h23de000b,32'hafdf000a,32'he7c10009,32'he7c00008,32'hafc20007,32'hc4610000,32'h20630003,32'h8fc30002,32'h46010000,32'h46020842,32'hc7c20003,32'hc4610000,32'h20230003,32'h46010000,32'h46020842,32'hc7c20004,32'hc4610000,32'h20230002,32'h46010002,32'hc7c10005,32'hc4600000,32'h20230001,32'h8fc10006,32'h143a004a,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0007,32'h23defff8,32'h0c0000ad,32'h23de0008,32'hafdf0007,32'h46030006,32'hafc20006,32'he7c00005,32'he7c10004,32'he7c20003,32'hafc30002,32'he7c30001,32'hafc10000,32'hc4830000,32'h20440000,32'h03e00008,32'h20010001,32'he4200000,32'h20410000,32'h46010002,32'hc4210000,32'h20210003,32'h8fc10000,32'hc4200000,32'h20210000,32'h8fc10001,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0002,32'h23defffd,32'h0c0000a4,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc30000,32'hc4200000,32'h20410000,32'h08000c1b,32'h8fc2000a,32'h8fc10002,32'hc7c20009,32'hc7c10007,32'hc7c00005,32'h08000bf6,32'h8fc2000a,32'h8fc10002,32'hc7c20009,32'hc7c10007,32'hc7c00005,32'h143a0007,32'h201a0002,32'h08000afa,32'h8fc3000a,32'h8fc10002,32'hc7c20009,32'hc7c10007,32'hc7c00005,32'h20220000,32'h8fdf000b,32'h23defff4,32'h0c00041e,32'h23de000c,32'hafdf000b,32'h8fc10001,32'h143a000e,32'h201a0001,32'h8fdf000b,32'h23defff4,32'h0c0003b7,32'h23de000c,32'hafdf000b,32'h20410000,32'hafc1000a,32'h8fc20002,32'h8c210000,32'h00220820,32'h8fc20000,32'h8fdf000a,32'h23defff5,32'h0c000421,32'h23de000b,32'hafdf000a,32'he7c00009,32'h8fc10001,32'h46000801,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003da,32'h23de000a,32'hafdf0009,32'he7c10008,32'he7c00007,32'h8fc10002,32'hc4210000,32'h20210002,32'h8fc10003,32'h46000801,32'hc7c10006,32'h8fdf0007,32'h23defff8,32'h0c0003d6,32'h23de0008,32'hafdf0007,32'h20410000,32'he7c10006,32'he7c00005,32'h8fc20002,32'hc4410000,32'h20220001,32'h8fc10003,32'h46000801,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0003d2,32'h23de0006,32'hafdf0005,32'h20810000,32'he7c00004,32'hafc30003,32'hafc40002,32'hafc20001,32'hafc10000,32'hc4a00000,32'h20650000,32'h8c840000,32'h00812020,32'h34840048,32'h3c040000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'he4200000,32'h20210000,32'h8fc10006,32'h46010002,32'hc4210000,32'h20210004,32'h8fc10005,32'h46000800,32'hc7c10007,32'h46000004,32'hc7c0000a,32'h08000c8e,32'he4200000,32'h20210000,32'h8fc10006,32'h46010002,32'hc4210000,32'h20210004,32'h8fc10005,32'h46000801,32'hc7c10007,32'h46000004,32'hc7c0000a,32'h143a000d,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c0003bd,32'h23de000c,32'hafdf000b,32'h8fc10001,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c00009b,32'h23de000c,32'hafdf000b,32'he7c0000a,32'h46010001,32'h46011042,32'hc7c20000,32'hc7c10009,32'h8fdf000a,32'h23defff5,32'h0c0000bb,32'h23de000b,32'hafdf000a,32'h46010006,32'he7c00009,32'hc7c10007,32'h46000006,32'hc7c00008,32'h08000c59,32'h46000801,32'hc7c10008,32'hc4200000,32'h34210030,32'h3c010000,32'h143a0007,32'h201a0003,32'h8fdf0009,32'h23defff6,32'h0c0003b7,32'h23de000a,32'hafdf0009,32'he7c00008,32'h8fc10001,32'h8fdf0008,32'h23defff7,32'h0c000947,32'h23de0009,32'hafdf0008,32'h46030046,32'h46010006,32'h46040086,32'h20610000,32'he7c00007,32'hafc20006,32'h8fc30001,32'h46020000,32'h46041082,32'hc7c40002,32'hc4620000,32'h20230003,32'h46020000,32'h46031082,32'hc7c30003,32'hc4620000,32'h20230002,32'h46010002,32'hc7c10004,32'hc4600000,32'h20230001,32'h8fc10005,32'h143a0064,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0006,32'h23defff9,32'h0c0000ad,32'h23de0007,32'hafdf0006,32'h46030006,32'hafc20005,32'he7c00004,32'he7c10003,32'he7c20002,32'hafc10001,32'he7c30000,32'hc4630000,32'h20430000,32'h03e00008,32'h20010001,32'he4200000,32'h20410000,32'h46010000,32'h46020842,32'hc7c20000,32'hc4210000,32'h20210003,32'h46010000,32'h46020842,32'hc7c20001,32'hc4610000,32'h20230002,32'h46010002,32'hc7c10002,32'hc4600000,32'h20230001,32'h8fc10003,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0004,32'h23defffb,32'h0c0000a4,32'h23de0005,32'hafdf0004,32'h46030006,32'hafc20003,32'he7c00002,32'he7c10001,32'he7c20000,32'hc4230000,32'h20410000,32'h03e00008,32'h20010001,32'he4200000,32'hc7c00005,32'h20410000,32'h03e00008,32'h20010002,32'he4200000,32'hc7c0000a,32'h20210000,32'h8fc10009,32'h03e00008,32'h20010003,32'he4200000,32'hc7c0000d,32'h20210000,32'h8fc10009,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h20010000,32'h08000be1,32'h20010001,32'h143a0003,32'h201a0000,32'h8fdf0010,32'h23deffef,32'h0c0000ad,32'h23de0011,32'hafdf0010,32'hc4200000,32'h20210005,32'h8fc10002,32'h08000be1,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0010,32'h23deffef,32'h0c000095,32'h23de0011,32'hafdf0010,32'hc7c0000f,32'h46000046,32'h8fdf0010,32'h23deffef,32'h0c0003c7,32'h23de0011,32'hafdf0010,32'he7c0000f,32'h8fc10003,32'h46000005,32'h46020000,32'hc7c20001,32'h46000802,32'hc7c1000d,32'hc4200000,32'h20210001,32'h8fc10006,32'h08000be1,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000f,32'h23defff0,32'h0c000095,32'h23de0010,32'hafdf000f,32'hc7c0000e,32'h46000046,32'h8fdf000f,32'h23defff0,32'h0c0003c3,32'h23de0010,32'hafdf000f,32'h20610000,32'he7c1000e,32'he7c0000d,32'h8fc30003,32'h46010045,32'h46020840,32'hc7c20000,32'h46010042,32'hc4610000,32'h20430000,32'h8fc20006,32'h46010002,32'hc4410000,32'h20220005,32'h46010001,32'hc7c10004,32'hc4400000,32'h20220004,32'h8fc10002,32'h143a0055,32'h201a0000,32'h20010000,32'h08000b95,32'h20010001,32'h143a0003,32'h201a0000,32'h8fdf000d,32'h23defff2,32'h0c0000ad,32'h23de000e,32'hafdf000d,32'hc4400000,32'h20220003,32'h8fc10002,32'h08000b95,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000d,32'h23defff2,32'h0c000095,32'h23de000e,32'hafdf000d,32'hc7c0000c,32'h46000046,32'h8fdf000d,32'h23defff2,32'h0c0003cb,32'h23de000e,32'hafdf000d,32'h20410000,32'he7c0000c,32'h8fc20003,32'h46000005,32'h46020000,32'hc7c20004,32'h46000802,32'hc7c1000a,32'hc4400000,32'h20220002,32'h8fc10006,32'h08000b95,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h0c000095,32'h23de000d,32'hafdf000c,32'hc7c0000b,32'h46000046,32'h8fdf000c,32'h23defff3,32'h0c0003c3,32'h23de000d,32'hafdf000c,32'h20810000,32'he7c2000b,32'he7c0000a,32'hafc20009,32'h8fc40003,32'h46020085,32'h46031080,32'hc7c30000,32'h46020082,32'hc4820000,32'h20640000,32'h8fc30006,32'h46020002,32'hc4620000,32'h20230003,32'h46010001,32'hc7c10001,32'hc4600000,32'h20230002,32'h8fc10002,32'h143a00a9,32'h201a0000,32'h344200c1,32'h3c020000,32'h20010000,32'h08000b45,32'h20010001,32'h143a0003,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c0000ad,32'h23de000a,32'hafdf0009,32'hc4400000,32'h20220001,32'h8fc10002,32'h08000b45,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0009,32'h23defff6,32'h0c000095,32'h23de000a,32'hafdf0009,32'hc7c00008,32'h46000046,32'h8fdf0009,32'h23defff6,32'h0c0003cb,32'h23de000a,32'hafdf0009,32'h20410000,32'he7c00008,32'h8fc20003,32'h46000005,32'h46020000,32'hc7c20004,32'h46000802,32'hc7c10005,32'hc4400000,32'h20220002,32'h8fc10006,32'h08000b45,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0008,32'h23defff7,32'h0c000095,32'h23de0009,32'hafdf0008,32'hc7c00007,32'h46000046,32'h8fdf0008,32'h23defff7,32'h0c0003c7,32'h23de0009,32'hafdf0008,32'he7c40007,32'hafc20006,32'he7c30005,32'he7c20004,32'hafc10003,32'hafc30002,32'he7c10001,32'he7c00000,32'h46040105,32'h46012100,32'h46041902,32'hc4840000,32'h20440001,32'h460418c2,32'hc4840000,32'h20640001,32'h460018c1,32'hc4830000,32'h20640000,32'h08000a30,32'h8fc20000,32'h8fc10001,32'hc7c20008,32'hc7c10006,32'hc7c00004,32'h08000914,32'h8fc20000,32'h8fc10001,32'hc7c20008,32'hc7c10006,32'hc7c00004,32'h143a0007,32'h201a0002,32'h080008df,32'h8fc20000,32'h8fc10001,32'hc7c20008,32'hc7c10006,32'hc7c00004,32'h143a0007,32'h201a0001,32'h8fdf0009,32'h23defff6,32'h0c0003b7,32'h23de000a,32'hafdf0009,32'he7c00008,32'h8fc10001,32'h46000801,32'hc7c10007,32'h8fdf0008,32'h23defff7,32'h0c0003da,32'h23de0009,32'hafdf0008,32'he7c10007,32'he7c00006,32'h8fc10001,32'hc4210000,32'h20210002,32'h8fc10002,32'h46000801,32'hc7c10005,32'h8fdf0006,32'h23defff9,32'h0c0003d6,32'h23de0007,32'hafdf0006,32'h20410000,32'he7c10005,32'he7c00004,32'h8fc20001,32'hc4410000,32'h20220001,32'h8fc10002,32'h46000801,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0003d2,32'h23de0005,32'hafdf0004,32'he7c00003,32'hafc30002,32'hafc10001,32'hafc20000,32'hc4800000,32'h20640000,32'h8c210000,32'h00810820,32'h34840048,32'h3c040000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'he4200000,32'h20210000,32'h8fc10006,32'h46010003,32'hc7c10005,32'h46010001,32'hc7c10007,32'h46000006,32'hc7c0000b,32'h08000aa6,32'h8fdf000c,32'h23defff3,32'h0c002471,32'h23de000d,32'hafdf000c,32'hc7c0000b,32'h143a0008,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h0c0003bd,32'h23de000d,32'hafdf000c,32'he7c0000b,32'h8fc10003,32'h46000004,32'hc7c0000a,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000b,32'h23defff4,32'h0c00009b,32'h23de000c,32'hafdf000b,32'he7c0000a,32'h46010001,32'h46011042,32'hc7c20005,32'hc7c10009,32'h8fdf000a,32'h23defff5,32'h0c0000bb,32'h23de000b,32'hafdf000a,32'h46010006,32'he7c00009,32'hc7c10007,32'h46000006,32'hc7c00008,32'h08000a7c,32'h46000801,32'hc7c10008,32'hc4200000,32'h34210030,32'h3c010000,32'h143a0007,32'h201a0003,32'h8fdf0009,32'h23defff6,32'h0c0003b7,32'h23de000a,32'hafdf0009,32'he7c00008,32'h8fc10003,32'h8fdf0008,32'h23defff7,32'h0c000947,32'h23de0009,32'hafdf0008,32'h46030086,32'h46020046,32'h46010006,32'he7c00007,32'h8fc10003,32'hc7c30000,32'hc7c20001,32'hc7c10002,32'h8fdf0007,32'h23defff8,32'h0c0009b8,32'h23de0008,32'hafdf0007,32'hafc20006,32'h8fc10003,32'hc7c50000,32'hc7c40001,32'hc7c30002,32'hc4220000,32'h20210002,32'hc4610000,32'h20230001,32'hc4600000,32'h20230000,32'h8fc10004,32'h143a0063,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0006,32'h23defff9,32'h0c0000ad,32'h23de0007,32'hafdf0006,32'he7c00005,32'h8fdf0005,32'h23defffa,32'h0c000947,32'h23de0006,32'hafdf0005,32'h46030006,32'h46040046,32'h46050086,32'hafc20004,32'hafc10003,32'he7c00002,32'he7c10001,32'he7c20000,32'hc4650000,32'h20430002,32'hc4640000,32'h20430001,32'hc4630000,32'h20430000,32'h03e00008,32'h46000800,32'hc7c1000c,32'h8fdf0012,32'h23deffed,32'h0c0000b6,32'h23de0013,32'hafdf0012,32'h46000800,32'hc7c10010,32'h46000802,32'hc7c10011,32'h8fdf0012,32'h23deffed,32'h0c0003fa,32'h23de0013,32'hafdf0012,32'he7c10011,32'he7c00010,32'h8fc10004,32'h46020840,32'h46021882,32'hc7c30006,32'hc7c20000,32'h46011042,32'hc7c20001,32'hc7c10005,32'h46000800,32'hc7c1000e,32'h46000802,32'hc7c1000f,32'h8fdf0010,32'h23deffef,32'h0c0003f6,32'h23de0011,32'hafdf0010,32'he7c1000f,32'he7c0000e,32'h8fc10004,32'h46040840,32'h46032102,32'hc7c40003,32'hc7c30000,32'h46011042,32'hc7c20001,32'hc7c10002,32'h46000802,32'hc7c1000d,32'h8fdf000e,32'h23defff1,32'h0c0003f2,32'h23de000f,32'hafdf000e,32'he7c2000d,32'h8fc10004,32'h46051080,32'h46032142,32'hc7c40006,32'hc7c30002,32'h46000882,32'hc7c10003,32'hc7c00005,32'h03e00008,32'h46000006,32'hc7c0000c,32'h143a0004,32'h201a0000,32'h8fdf000d,32'h23defff2,32'h0c0003c0,32'h23de000e,32'hafdf000d,32'he7c0000c,32'h8fc10004,32'h46000800,32'hc7c1000a,32'h46000802,32'hc7c1000b,32'h8fdf000c,32'h23defff3,32'h0c0003cb,32'h23de000d,32'hafdf000c,32'he7c3000b,32'he7c0000a,32'h8fc10004,32'h460110c2,32'hc7c20003,32'hc7c10002,32'h46000800,32'hc7c10008,32'h46000802,32'hc7c10009,32'h8fdf000a,32'h23defff5,32'h0c0003c7,32'h23de000b,32'hafdf000a,32'he7c30009,32'he7c00008,32'h8fc10004,32'h460110c2,32'hc7c20006,32'hc7c10005,32'h46000802,32'hc7c10007,32'h8fdf0008,32'h23defff7,32'h0c0003c3,32'h23de0009,32'hafdf0008,32'he7c60007,32'he7c10006,32'he7c40005,32'hafc10004,32'he7c20003,32'he7c50002,32'he7c00001,32'he7c30000,32'h46030182,32'h03e00008,32'h46000800,32'hc7c1000d,32'h46000802,32'hc7c1000e,32'h8fdf000f,32'h23defff0,32'h0c0003fa,32'h23de0010,32'hafdf000f,32'he7c1000e,32'he7c0000d,32'h8fc10002,32'h46011042,32'hc7c20000,32'hc7c10003,32'h46000800,32'hc7c1000b,32'h46000802,32'hc7c1000c,32'h8fdf000d,32'h23defff2,32'h0c0003f6,32'h23de000e,32'hafdf000d,32'he7c2000c,32'he7c0000b,32'h8fc10002,32'h46011082,32'hc7c20001,32'hc7c10000,32'h46000800,32'hc7c10009,32'h46000802,32'hc7c1000a,32'h8fdf000b,32'h23defff4,32'h0c0003f2,32'h23de000c,32'hafdf000b,32'he7c2000a,32'h8fc10002,32'h46000882,32'hc7c10003,32'hc7c00001,32'h03e00008,32'h46000006,32'hc7c00009,32'h143a0004,32'h201a0000,32'h8fdf000a,32'h23defff5,32'h0c0003c0,32'h23de000b,32'hafdf000a,32'he7c00009,32'h8fc10002,32'h46000800,32'hc7c10007,32'h46000802,32'hc7c10008,32'h8fdf0009,32'h23defff6,32'h0c0003cb,32'h23de000a,32'hafdf0009,32'he7c00008,32'h8fc10002,32'h8fdf0008,32'h23defff7,32'h0c0000bb,32'h23de0009,32'hafdf0008,32'h46010006,32'he7c00007,32'hc7c10001,32'h46000800,32'hc7c10005,32'h46000802,32'hc7c10006,32'h8fdf0007,32'h23defff8,32'h0c0003c7,32'h23de0008,32'hafdf0007,32'he7c00006,32'h8fc10002,32'h8fdf0006,32'h23defff9,32'h0c0000bb,32'h23de0007,32'hafdf0006,32'h46010006,32'he7c00005,32'hc7c10003,32'h46000802,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0003c3,32'h23de0006,32'hafdf0005,32'he7c00004,32'h8fc10002,32'h8fdf0004,32'h23defffb,32'h0c0000bb,32'h23de0005,32'hafdf0004,32'he7c10003,32'hafc10002,32'he7c20001,32'he7c00000,32'h03e00008,32'h20010001,32'he4200000,32'h20210000,32'h8fc10006,32'h46010003,32'hc7c10005,32'h8fdf0007,32'h23defff8,32'h0c002471,32'h23de0008,32'hafdf0007,32'h8fdf0007,32'h23defff8,32'h0c00034a,32'h23de0008,32'hafdf0007,32'hafc20006,32'h8fc10004,32'hc7c20000,32'hc7c10001,32'hc7c00002,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0006,32'h23defff9,32'h0c00009b,32'h23de0007,32'hafdf0006,32'he7c00005,32'h8fdf0005,32'h23defffa,32'h0c000338,32'h23de0006,32'hafdf0005,32'hafc20004,32'h8fc10003,32'h20220000,32'h8fdf0004,32'h23defffb,32'h0c0003cf,32'h23de0005,32'hafdf0004,32'hafc20003,32'he7c00002,32'he7c10001,32'he7c20000,32'h03e00008,32'h20010001,32'h03e00008,32'h20010002,32'h03e00008,32'h20010003,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c000867,32'h23de0006,32'hafdf0005,32'h8fc20003,32'h8fc10004,32'hc7c20002,32'hc7c10000,32'hc7c00001,32'h20050001,32'h20040000,32'h20030002,32'h143a0014,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c000867,32'h23de0006,32'hafdf0005,32'h8fc20003,32'h8fc10004,32'hc7c20000,32'hc7c10001,32'hc7c00002,32'h20050000,32'h20040002,32'h20030001,32'h143a0025,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c000867,32'h23de0006,32'hafdf0005,32'hafc10004,32'hafc20003,32'he7c10002,32'he7c20001,32'he7c00000,32'h20050002,32'h20040001,32'h20030000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'he4200000,32'hc7c0000b,32'h20210000,32'h8fc10008,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h0c000095,32'h23de000d,32'hafdf000c,32'h46020046,32'hc4220000,32'h00410820,32'h8fc20009,32'h46000005,32'h46020000,32'hc7c20000,32'h46000802,32'hc7c1000b,32'hc4400000,32'h00411020,32'h8fc20006,32'h8fc10001,32'h03e00008,32'h20010000,32'h143a0003,32'h201a0000,32'h8fdf000c,32'h23defff3,32'h0c000095,32'h23de000d,32'hafdf000c,32'h46020046,32'h46010006,32'he7c0000b,32'hc4220000,32'h00610820,32'h8fc30009,32'h46010045,32'h46020840,32'hc7c20002,32'h46010042,32'hc4610000,32'h00411820,32'h8fc10003,32'h46010003,32'hc4210000,32'h00410820,32'h8fc20006,32'h8fc10005,32'h46010001,32'hc7c10004,32'h8fdf000b,32'h23defff4,32'h0c0002bf,32'h23de000c,32'hafdf000b,32'hc4800000,32'h00622020,32'h8fc30009,32'h8fc20005,32'h8fdf000b,32'h23defff4,32'h0c000299,32'h23de000c,32'hafdf000b,32'h8fc1000a,32'h20220000,32'h8fdf000b,32'h23defff4,32'h0c0000a4,32'h23de000c,32'hafdf000b,32'hafc1000a,32'hc4800000,32'h00622020,32'h8fc30006,32'h8fc20005,32'h8fdf000a,32'h23defff5,32'h0c0003bd,32'h23de000b,32'hafdf000a,32'h20410000,32'hafc10009,32'h8fc20007,32'h8fdf0009,32'h23defff6,32'h0c0003cf,32'h23de000a,32'hafdf0009,32'hafc20008,32'h8fc10007,32'h143a0063,32'h201a0000,32'h344200c1,32'h3c020000,32'h8fdf0008,32'h23defff7,32'h0c0000ad,32'h23de0009,32'hafdf0008,32'h46030006,32'hafc10007,32'hafc20006,32'hafc30005,32'he7c00004,32'hafc40003,32'he7c10002,32'hafc50001,32'he7c20000,32'hc4c30000,32'h00433020,32'h03e00008,32'hac410000,32'h20420000,32'h8fc20000,32'h8fdf0001,32'h23defffe,32'h0c000813,32'h23de0002,32'hafdf0001,32'h20010000,32'h8fdf0001,32'h23defffe,32'h0c000832,32'h23de0002,32'hafdf0001,32'h20010000,32'h8fdf0001,32'h23defffe,32'h0c0007f6,32'h23de0002,32'hafdf0001,32'h8fdf0001,32'h23defffe,32'h0c0004e5,32'h23de0002,32'hafdf0001,32'h8fdf0001,32'h23defffe,32'h0c000432,32'h23de0002,32'hafdf0001,32'hafc10000,32'h8f610001,32'h08000832,32'h20410001,32'hac610000,32'h00621820,32'h8fc20000,32'h03e00008,32'h145a0002,32'h201affff,32'h3463008f,32'h3c030000,32'h8c420000,32'h20220000,32'h8fdf0001,32'h23defffe,32'h0c0007f8,32'h23de0002,32'hafdf0001,32'h20410000,32'hafc10000,32'h20020000,32'h03e00008,32'h00010820,32'hac430000,32'h8fc30001,32'h00221020,32'h8fc20000,32'h8fdf0002,32'h23defffd,32'h0c000813,32'h23de0003,32'hafdf0002,32'h20610000,32'hafc20001,32'h20230001,32'h8fc10000,32'h08002461,32'h20210001,32'h8fc10000,32'h143a0004,32'h201affff,32'h8c210000,32'h20410000,32'h20220000,32'h8fdf0001,32'h23defffe,32'h0c0007f8,32'h23de0002,32'hafdf0001,32'h20410000,32'hafc10000,32'h20020000,32'h03e00008,32'h00010820,32'hac430000,32'h8fc30001,32'h00221020,32'h8fc20000,32'h8fdf0002,32'h23defffd,32'h0c0007f8,32'h23de0003,32'hafdf0002,32'h20610000,32'hafc10001,32'h20430001,32'h8fc20000,32'h08002461,32'h2002ffff,32'h20210001,32'h8fc10000,32'h143a0005,32'h201affff,32'h8fdf0001,32'h23defffe,32'h0c002473,32'h23de0002,32'hafdf0001,32'hafc10000,32'h080007df,32'h20010000,32'h080007df,32'h20210001,32'h8fc10000,32'h03e00008,32'hac220000,32'h8fc20000,32'h20210000,32'h8fc10001,32'h143a0006,32'h201a0000,32'h8fdf0002,32'h23defffd,32'h0c000649,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc10000,32'h03e00008,32'h13800002,32'h0341e02a,32'h201a003c,32'h34420047,32'h3c020000,32'h03e00008,32'h20010001,32'h8fdf0013,32'h23deffec,32'h0c000538,32'h23de0014,32'hafdf0013,32'h8fc2000b,32'h8fc10006,32'h080007dd,32'h143a0002,32'h201a0000,32'h8fc10005,32'h080007d2,32'h8fdf0013,32'h23deffec,32'h0c0002eb,32'h23de0014,32'hafdf0013,32'h20610000,32'h20020000,32'h080007cb,32'h20020001,32'h145a0003,32'h201a0000,32'h8fc20008,32'h14ba000e,32'h201a0002,32'h080007d2,32'he4400000,32'h20220002,32'h8fc10006,32'hc4200000,32'h34210032,32'h3c010000,32'h080007bf,32'h46000803,32'hc7c10012,32'h8fdf0013,32'h23deffec,32'h0c0000bb,32'h23de0014,32'hafdf0013,32'h46010006,32'he7c00012,32'hc7c10011,32'h8fdf0012,32'h23deffed,32'h0c0002a3,32'h23de0013,32'hafdf0012,32'hc7c00011,32'h143a0012,32'h201a0000,32'h8fdf0012,32'h23deffed,32'h0c0000ad,32'h23de0013,32'hafdf0012,32'he7c00011,32'hc4400000,32'h20220002,32'he4400000,32'h20220001,32'h8fc10006,32'hc4200000,32'h34210032,32'h3c010000,32'h0800079e,32'h46000803,32'hc7c10010,32'h8fdf0011,32'h23deffee,32'h0c0000bb,32'h23de0012,32'hafdf0011,32'h46010006,32'he7c00010,32'hc7c1000f,32'h8fdf0010,32'h23deffef,32'h0c0002a3,32'h23de0011,32'hafdf0010,32'hc7c0000f,32'h143a0012,32'h201a0000,32'h8fdf0010,32'h23deffef,32'h0c0000ad,32'h23de0011,32'hafdf0010,32'he7c0000f,32'hc4400000,32'h20220001,32'he4400000,32'h20220000,32'h8fc10006,32'hc4200000,32'h34210032,32'h3c010000,32'h0800077d,32'h46000803,32'hc7c1000e,32'h8fdf000f,32'h23defff0,32'h0c0000bb,32'h23de0010,32'hafdf000f,32'h46010006,32'he7c0000e,32'hc7c1000d,32'h8fdf000e,32'h23defff1,32'h0c0002a3,32'h23de000f,32'hafdf000e,32'hc7c0000d,32'h143a0012,32'h201a0000,32'h8fdf000e,32'h23defff1,32'h0c0000ad,32'h23de000f,32'hafdf000e,32'he7c0000d,32'hc4400000,32'h20620000,32'h14ba0065,32'h201a0003,32'hacc20000,32'h00e63020,32'h8fc70001,32'h8fc60000,32'h20420000,32'hac460000,32'h8fc60002,32'hac450001,32'h8fc50003,32'hac450002,32'h8fc50004,32'hac440003,32'h8fc40005,32'hac430004,32'h8fc30006,32'hac430005,32'h8fc30007,32'hac430006,32'h8fc3000c,32'hac430007,32'h8fc30009,32'hac430008,32'h8fc3000a,32'hac410009,32'h8fc1000b,32'hac41000a,32'h23bd000b,32'h23a20000,32'h8fdf000d,32'h23defff2,32'h0c002469,32'h23de000e,32'hafdf000d,32'h20810000,32'hafc1000b,32'hafc3000c,32'hc4a00000,32'h34a50032,32'h3c050000,32'h20040004,32'h00031820,32'h8fc30008,32'h08000735,32'h20030001,32'h145a0003,32'h201a0002,32'h8fc20003,32'he4400000,32'h20220002,32'h8fc1000b,32'h8fdf000c,32'h23defff3,32'h0c00042d,32'h23de000d,32'hafdf000c,32'h8fdf000c,32'h23defff3,32'h0c002482,32'h23de000d,32'hafdf000c,32'he4400000,32'h20220001,32'h8fc1000b,32'h8fdf000c,32'h23defff3,32'h0c00042d,32'h23de000d,32'hafdf000c,32'h8fdf000c,32'h23defff3,32'h0c002482,32'h23de000d,32'hafdf000c,32'he4400000,32'h20220000,32'h8fc1000b,32'h8fdf000c,32'h23defff3,32'h0c00042d,32'h23de000d,32'hafdf000c,32'h8fdf000c,32'h23defff3,32'h0c002482,32'h23de000d,32'hafdf000c,32'hafc1000b,32'h0800072e,32'h145a0002,32'h201a0000,32'h8fc20005,32'h8fdf000b,32'h23defff4,32'h0c002469,32'h23de000c,32'hafdf000b,32'h20410000,32'hc4600000,32'h34630032,32'h3c030000,32'h20020003,32'he4400000,32'h20220002,32'h8fc1000a,32'h8fdf000b,32'h23defff4,32'h0c002482,32'h23de000c,32'hafdf000b,32'he4400000,32'h20220001,32'h8fc1000a,32'h8fdf000b,32'h23defff4,32'h0c002482,32'h23de000c,32'hafdf000b,32'he4400000,32'h20220000,32'h8fc1000a,32'h8fdf000b,32'h23defff4,32'h0c002482,32'h23de000c,32'hafdf000b,32'hafc1000a,32'h8fdf000a,32'h23defff5,32'h0c002469,32'h23de000b,32'hafdf000a,32'h20410000,32'hc4600000,32'h34630032,32'h3c030000,32'h20020003,32'he4400000,32'h20220001,32'h8fc10009,32'h8fdf000a,32'h23defff5,32'h0c002482,32'h23de000b,32'hafdf000a,32'he4400000,32'h20220000,32'h8fc10009,32'h8fdf000a,32'h23defff5,32'h0c002482,32'h23de000b,32'hafdf000a,32'hafc10009,32'h8fdf0009,32'h23defff6,32'h0c002469,32'h23de000a,32'hafdf0009,32'h20410000,32'hafc10008,32'hc4600000,32'h34630032,32'h3c030000,32'h20020002,32'h8fdf0008,32'h23defff7,32'h0c0000a4,32'h23de0009,32'hafdf0008,32'h8fdf0008,32'h23defff7,32'h0c002482,32'h23de0009,32'hafdf0008,32'he4400000,32'h20220002,32'h8fc10007,32'h8fdf0008,32'h23defff7,32'h0c002482,32'h23de0009,32'hafdf0008,32'he4400000,32'h20220001,32'h8fc10007,32'h8fdf0008,32'h23defff7,32'h0c002482,32'h23de0009,32'hafdf0008,32'he4400000,32'h20220000,32'h8fc10007,32'h8fdf0008,32'h23defff7,32'h0c002482,32'h23de0009,32'hafdf0008,32'hafc10007,32'h8fdf0007,32'h23defff8,32'h0c002469,32'h23de0008,32'hafdf0007,32'h20410000,32'hc4600000,32'h34630032,32'h3c030000,32'h20020003,32'he4400000,32'h20220002,32'h8fc10006,32'h8fdf0007,32'h23defff8,32'h0c002482,32'h23de0008,32'hafdf0007,32'he4400000,32'h20220001,32'h8fc10006,32'h8fdf0007,32'h23defff8,32'h0c002482,32'h23de0008,32'hafdf0007,32'he4400000,32'h20220000,32'h8fc10006,32'h8fdf0007,32'h23defff8,32'h0c002482,32'h23de0008,32'hafdf0007,32'hafc10006,32'h8fdf0006,32'h23defff9,32'h0c002469,32'h23de0007,32'hafdf0006,32'h20410000,32'hafc10005,32'hc4600000,32'h34630032,32'h3c030000,32'h20020003,32'h8fdf0005,32'h23defffa,32'h0c002473,32'h23de0006,32'hafdf0005,32'hafc10004,32'h8fdf0004,32'h23defffb,32'h0c002473,32'h23de0005,32'hafdf0004,32'hafc10003,32'h8fdf0003,32'h23defffc,32'h0c002473,32'h23de0004,32'hafdf0003,32'hafc10002,32'hafc20001,32'h03e00008,32'h20010000,32'h143a0003,32'h201affff,32'h34420048,32'h3c020000,32'h8fdf0001,32'h23defffe,32'h0c002473,32'h23de0002,32'hafdf0001,32'hafc10000,32'h03e00008,32'he4200000,32'h20210002,32'h46010002,32'h46011040,32'h46080842,32'h46090842,32'h46031080,32'h460618c2,32'h460a38c2,32'h46021882,32'h460418c2,32'hc4400000,32'h34420017,32'h3c020000,32'he4400000,32'h20220001,32'h46050002,32'h460b2940,32'h460b62c2,32'h46090b02,32'hc7c90011,32'h46092940,32'h46096242,32'h460a3b02,32'hc7ca000b,32'h46055142,32'h46041a82,32'hc7c4000c,32'hc4400000,32'h34420017,32'h3c020000,32'he4400000,32'h20220000,32'h8fc10001,32'h46040002,32'h460a2100,32'h460b5282,32'hc7cb000d,32'h46080a82,32'hc7c8000e,32'h46082100,32'h46094202,32'hc7c90007,32'h46063a02,32'hc7c70012,32'hc7c60009,32'h46052102,32'hc7c50008,32'h46021902,32'hc7c3000f,32'hc7c2000a,32'hc4200000,32'h34210017,32'h3c010000,32'he4200000,32'h20210002,32'h8fc10000,32'h46001000,32'hc7c20018,32'h46000802,32'hc7c10010,32'h8fdf0019,32'h23deffe6,32'h0c0000bb,32'h23de001a,32'hafdf0019,32'h46020006,32'he7c00018,32'hc7c2000d,32'h46001000,32'hc7c20017,32'h46000802,32'hc7c10012,32'h8fdf0018,32'h23deffe7,32'h0c0000bb,32'h23de0019,32'hafdf0018,32'h46020006,32'he7c00017,32'hc7c20007,32'h46000802,32'hc7c1000f,32'h8fdf0017,32'h23deffe8,32'h0c0000bb,32'h23de0018,32'hafdf0017,32'hc7c00008,32'he4400000,32'h20220001,32'h8fc10000,32'h46001000,32'hc7c20016,32'h46000802,32'hc7c10010,32'h8fdf0017,32'h23deffe8,32'h0c0000bb,32'h23de0018,32'hafdf0017,32'h46020006,32'he7c00016,32'hc7c2000e,32'h46001000,32'hc7c20015,32'h46000802,32'hc7c10012,32'h8fdf0016,32'h23deffe9,32'h0c0000bb,32'h23de0017,32'hafdf0016,32'h46020006,32'he7c00015,32'hc7c20009,32'h46000802,32'hc7c1000f,32'h8fdf0015,32'h23deffea,32'h0c0000bb,32'h23de0016,32'hafdf0015,32'hc7c0000a,32'he4400000,32'h20220000,32'h8fc10000,32'h46001000,32'hc7c20014,32'h46000802,32'hc7c10010,32'h8fdf0015,32'h23deffea,32'h0c0000bb,32'h23de0016,32'hafdf0015,32'h46020006,32'he7c00014,32'hc7c20011,32'h46001000,32'hc7c20013,32'h46000802,32'hc7c10012,32'h8fdf0014,32'h23deffeb,32'h0c0000bb,32'h23de0015,32'hafdf0014,32'h46020006,32'he7c00013,32'hc7c2000b,32'h46000802,32'hc7c1000f,32'h8fdf0013,32'h23deffec,32'h0c0000bb,32'h23de0014,32'hafdf0013,32'h46060006,32'he7c40012,32'he7c00011,32'he7c50010,32'he7c3000f,32'he7c2000e,32'he7c1000d,32'hc7c6000c,32'hc4450000,32'h20220002,32'hc4440000,32'h20220001,32'hc4430000,32'h20220000,32'h8fc10000,32'h46011842,32'hc7c30002,32'h46011082,32'hc7c20003,32'hc7c10004,32'h8fdf000d,32'h23defff2,32'h0c002471,32'h23de000e,32'hafdf000d,32'h46040006,32'he7c3000c,32'he7c9000b,32'he7c6000a,32'he7ca0009,32'he7c80008,32'he7c00007,32'h46010001,32'h46012842,32'h46005802,32'h46043ac2,32'h460b5280,32'h46013ac2,32'h46005282,32'h46042a82,32'h46001242,32'h46094200,32'h46002a42,32'h46014202,32'h46043a02,32'h46083181,32'h46003a02,32'hc7c70002,32'h46013182,32'h46042982,32'hc7c50003,32'hc7c40005,32'h460110c2,32'hc7c20004,32'hc7c10006,32'h8fdf0007,32'h23defff8,32'h0c00016d,32'h23de0008,32'hafdf0007,32'h46010006,32'he7c00006,32'hc4410000,32'h20220002,32'h8fc10001,32'h8fdf0006,32'h23defff9,32'h0c0000e6,32'h23de0007,32'hafdf0006,32'h46010006,32'he7c00005,32'hc4410000,32'h20220002,32'h8fc10001,32'h8fdf0005,32'h23defffa,32'h0c00016d,32'h23de0006,32'hafdf0005,32'h46010006,32'he7c00004,32'hc4410000,32'h20220001,32'h8fc10001,32'h8fdf0004,32'h23defffb,32'h0c0000e6,32'h23de0005,32'hafdf0004,32'h46010006,32'he7c00003,32'hc4410000,32'h20220001,32'h8fc10001,32'h8fdf0003,32'h23defffc,32'h0c00016d,32'h23de0004,32'hafdf0003,32'h46010006,32'he7c00002,32'hc4410000,32'h20220000,32'h8fc10001,32'h8fdf0002,32'h23defffd,32'h0c0000e6,32'h23de0003,32'hafdf0002,32'hafc20001,32'hafc10000,32'hc4600000,32'h20430000,32'h03e00008,32'he4200000,32'h20210000,32'h3421008d,32'h3c010000,32'h8fdf0004,32'h23defffb,32'h0c002482,32'h23de0005,32'hafdf0004,32'he4200000,32'h20210002,32'h8fc10001,32'h46000802,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0000e6,32'h23de0005,32'hafdf0004,32'hc7c00002,32'he4400000,32'h20220000,32'h8fc10001,32'h46000802,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c00016d,32'h23de0005,32'hafdf0004,32'h46010006,32'he7c00003,32'hc7c10002,32'h8fdf0003,32'h23defffc,32'h0c0000e6,32'h23de0004,32'hafdf0003,32'h46010006,32'he7c00002,32'hc7c10000,32'h8fdf0002,32'h23defffd,32'h0c00042d,32'h23de0003,32'hafdf0002,32'h8fdf0002,32'h23defffd,32'h0c002482,32'h23de0003,32'hafdf0002,32'hafc10001,32'he4400000,32'h20220001,32'h3421008a,32'h3c010000,32'h8fdf0001,32'h23defffe,32'h0c002471,32'h23de0002,32'hafdf0001,32'h8fdf0001,32'h23defffe,32'h0c00016d,32'h23de0002,32'hafdf0001,32'he7c00000,32'h8fdf0000,32'h23deffff,32'h0c00042d,32'h23de0001,32'hafdf0000,32'h8fdf0000,32'h23deffff,32'h0c002482,32'h23de0001,32'hafdf0000,32'h8fdf0000,32'h23deffff,32'h0c002473,32'h23de0001,32'hafdf0000,32'h03e00008,32'he4200000,32'h20610002,32'h46010001,32'hc4210000,32'h20410002,32'hc4200000,32'h20210002,32'he4800000,32'h20640001,32'h46010001,32'hc4810000,32'h20440001,32'hc4800000,32'h20240001,32'he4800000,32'h20640000,32'h34630087,32'h3c030000,32'h46010001,32'hc4610000,32'h20430000,32'h8fc20006,32'hc4400000,32'h20220000,32'h8fc10000,32'he4200000,32'h20210002,32'h8fc10009,32'h46010002,32'hc7c10005,32'h8fdf000a,32'h23defff5,32'h0c002471,32'h23de000b,32'hafdf000a,32'hc7c00003,32'he4400000,32'h20220001,32'h8fc10009,32'h8fdf000a,32'h23defff5,32'h0c002471,32'h23de000b,32'hafdf000a,32'hafc10009,32'hc7c00002,32'he4400000,32'h20220000,32'h342100e2,32'h3c010000,32'h46010002,32'hc7c10007,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'hc7c00003,32'he4200000,32'h20210002,32'h8fc10008,32'h8fdf0009,32'h23defff6,32'h0c002471,32'h23de000a,32'hafdf0009,32'hafc20008,32'he7c00007,32'hafc10006,32'he4640000,32'h20430001,32'hc4640000,32'h34630032,32'h3c030000,32'he4620000,32'h20430000,32'h344200df,32'h3c020000,32'he4440000,32'h20220002,32'h46052102,32'hc4450000,32'h34420019,32'h3c020000,32'h46020902,32'hc7c20005,32'he4420000,32'h20220001,32'h46021882,32'hc7c30003,32'hc4420000,32'h34420018,32'h3c020000,32'he4420000,32'h20220000,32'h342100e5,32'h3c010000,32'h46031082,32'hc4230000,32'h34210019,32'h3c010000,32'h46000882,32'hc7c10002,32'h8fdf0006,32'h23defff9,32'h0c00016d,32'h23de0007,32'hafdf0006,32'h46010006,32'he7c00005,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0000e6,32'h23de0006,32'hafdf0005,32'he7c00004,32'h8fdf0004,32'h23defffb,32'h0c00042d,32'h23de0005,32'hafdf0004,32'h8fdf0004,32'h23defffb,32'h0c002482,32'h23de0005,32'hafdf0004,32'he7c00003,32'h8fdf0003,32'h23defffc,32'h0c00016d,32'h23de0004,32'hafdf0003,32'h46010006,32'he7c00002,32'hc7c10001,32'h8fdf0002,32'h23defffd,32'h0c0000e6,32'h23de0003,32'hafdf0002,32'he7c00001,32'h8fdf0001,32'h23defffe,32'h0c00042d,32'h23de0002,32'hafdf0001,32'h8fdf0001,32'h23defffe,32'h0c002482,32'h23de0002,32'hafdf0001,32'he4400000,32'h20220002,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c002482,32'h23de0002,32'hafdf0001,32'he4400000,32'h20220001,32'h8fc10000,32'h8fdf0001,32'h23defffe,32'h0c002482,32'h23de0002,32'hafdf0001,32'hafc10000,32'he4400000,32'h20220000,32'h34210084,32'h3c010000,32'h8fdf0000,32'h23deffff,32'h0c002482,32'h23de0001,32'hafdf0000,32'h03e00008,32'h46010002,32'hc4210000,32'h3421001a,32'h3c010000,32'h03e00008,32'h46000006,32'hc4200002,32'h03e00008,32'h00010820,32'h8c210001,32'h03e00008,32'h00010820,32'h8c210000,32'h03e00008,32'h00010820,32'h8c210001,32'h03e00008,32'h00010820,32'h8c210000,32'h03e00008,32'h00010820,32'h8c210007,32'h03e00008,32'hac220000,32'h20210000,32'h8c210006,32'h03e00008,32'h8c210000,32'h20210000,32'h8c210006,32'h03e00008,32'h00010820,32'h8c210005,32'h03e00008,32'h00010820,32'h8c210004,32'h03e00008,32'h00010820,32'h8c210003,32'h03e00008,32'h00010820,32'h8c210002,32'h03e00008,32'h00010820,32'h8c210001,32'h03e00008,32'h00010820,32'h8c210000,32'h03e00008,32'h00010820,32'h8c21000a,32'h03e00008,32'hc4200000,32'h20210002,32'h8c210009,32'h03e00008,32'hc4200000,32'h20210001,32'h8c210009,32'h03e00008,32'hc4200000,32'h20210000,32'h8c210009,32'h03e00008,32'hc4200000,32'h20210002,32'h8c210008,32'h03e00008,32'hc4200000,32'h20210001,32'h8c210008,32'h03e00008,32'hc4200000,32'h20210000,32'h8c210008,32'h03e00008,32'hc4200000,32'h20210001,32'h8c210007,32'h03e00008,32'hc4200000,32'h20210000,32'h8c210007,32'h03e00008,32'hc4200000,32'h20210002,32'h8c210005,32'h03e00008,32'hc4200000,32'h20210001,32'h8c210005,32'h03e00008,32'hc4200000,32'h20210000,32'h8c210005,32'h03e00008,32'h00010820,32'h8c210004,32'h03e00008,32'hc4200000,32'h20210002,32'h8c210004,32'h03e00008,32'hc4200000,32'h20210001,32'h8c210004,32'h03e00008,32'hc4200000,32'h20210000,32'h8c210004,32'h03e00008,32'h00010820,32'h8c210003,32'h03e00008,32'h00010820,32'h8c210006,32'h03e00008,32'h00010820,32'h8c210002,32'h03e00008,32'h00010820,32'h8c210001,32'h03e00008,32'h00010820,32'h8c210000,32'h03e00008,32'he4200000,32'h20210002,32'h46010000,32'h46020842,32'hc4420000,32'h20620002,32'hc4410000,32'h20420002,32'hc4800000,32'h20240002,32'he4800000,32'h20240001,32'h46010000,32'h46020842,32'hc4820000,32'h20640001,32'hc4810000,32'h20440001,32'hc4800000,32'h20240001,32'he4800000,32'h20240000,32'h46010000,32'h46020842,32'hc4820000,32'h20640000,32'hc4810000,32'h20440000,32'hc4800000,32'h20240000,32'h03e00008,32'he4200000,32'h20210002,32'h46000802,32'hc4410000,32'h20220002,32'he4410000,32'h20220001,32'h46000842,32'hc4410000,32'h20220001,32'he4410000,32'h20220000,32'h46000842,32'hc4410000,32'h20220000,32'h03e00008,32'he4200000,32'h20210002,32'h46010000,32'hc4410000,32'h20420002,32'hc4600000,32'h20230002,32'he4600000,32'h20230001,32'h46010000,32'hc4610000,32'h20430001,32'hc4600000,32'h20230001,32'he4600000,32'h20230000,32'h46010000,32'hc4610000,32'h20430000,32'hc4600000,32'h20230000,32'h03e00008,32'he4200000,32'h20210002,32'h46000800,32'h46020002,32'hc4420000,32'h20420002,32'hc4610000,32'h20230002,32'he4610000,32'h20230001,32'h46020840,32'h46020082,32'hc4620000,32'h20430001,32'hc4610000,32'h20230001,32'he4610000,32'h20230000,32'h46020840,32'h46020082,32'hc4620000,32'h20430000,32'hc4610000,32'h20230000,32'h03e00008,32'h46010000,32'h46020842,32'hc4210000,32'h20210002,32'h46010000,32'h46011842,32'hc4430000,32'h20220001,32'h46001802,32'hc4430000,32'h20220000,32'h03e00008,32'h46010000,32'h46020842,32'hc4220000,32'h20410002,32'hc4210000,32'h20210002,32'h46010000,32'h46020842,32'hc4620000,32'h20430001,32'hc4610000,32'h20230001,32'h46010002,32'hc4610000,32'h20430000,32'hc4600000,32'h20230000,32'h03e00008,32'he4200000,32'h20210002,32'h46000802,32'hc4410000,32'h20220002,32'he4410000,32'h20220001,32'h46000842,32'hc4410000,32'h20220001,32'he4410000,32'h20220000,32'h46000842,32'hc4410000,32'h20220000,32'h8fc10001,32'hc4200000,32'h34210030,32'h3c010000,32'h08000327,32'h46010003,32'hc7c10004,32'hc4200000,32'h3421001b,32'h3c010000,32'h08000323,32'h46010003,32'hc7c10004,32'hc4200000,32'h34210030,32'h3c010000,32'h143a0007,32'h201a0000,32'h8fc10000,32'h143a0010,32'h201a0000,32'h8fdf0005,32'h23defffa,32'h0c0000ad,32'h23de0006,32'hafdf0005,32'he7c00004,32'h46000004,32'h46000800,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0000bb,32'h23de0005,32'hafdf0004,32'h46010006,32'he7c00003,32'hc4410000,32'h20220002,32'h8fc10001,32'h46000800,32'hc7c10002,32'h8fdf0003,32'h23defffc,32'h0c0000bb,32'h23de0004,32'hafdf0003,32'h46010006,32'he7c00002,32'hc4410000,32'h20220001,32'h8fc10001,32'h8fdf0002,32'h23defffd,32'h0c0000bb,32'h23de0003,32'hafdf0002,32'hafc10001,32'hafc20000,32'hc4600000,32'h20230000,32'h03e00008,32'he4200000,32'h20210002,32'hc4400000,32'h20420002,32'he4600000,32'h20230001,32'hc4600000,32'h20430001,32'he4600000,32'h20230000,32'hc4600000,32'h20430000,32'h080002d3,32'hc4400000,32'h34420032,32'h3c020000,32'h03e00008,32'he4200000,32'h20210002,32'he4400000,32'h20220001,32'he4400000,32'h20220000,32'h03e00008,32'he4220000,32'h20210002,32'he4410000,32'h20220001,32'he4400000,32'h20220000,32'h03e00008,32'h00010820,32'h03e00008,32'h2021fffb,32'h13800003,32'h0341e02a,32'h201a0005,32'h00220820,32'h03e00008,32'h46000006,32'h08002471,32'h143a0002,32'h201a0000,32'h03e00008,32'hc4200000,32'h34210032,32'h3c010000,32'h03e00008,32'hc4200000,32'h34210030,32'h3c010000,32'h03e00008,32'hc4200000,32'h3421001b,32'h3c010000,32'h143a0005,32'h201a0000,32'h8fdf0001,32'h23defffe,32'h0c00009b,32'h23de0002,32'hafdf0001,32'hc7c00000,32'h143a0011,32'h201a0000,32'h8fdf0001,32'h23defffe,32'h0c0000ad,32'h23de0002,32'hafdf0001,32'he7c00000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'h145a0003,32'h201a0000,32'h03e00008,32'h00020820,32'h143a0003,32'h201a0000,32'h03e00008,32'hc0200000,32'he0010000,32'h46010001,32'hc4210000,32'h34210031,32'h3c010000,32'h080001ff,32'h03e00008,32'h46000800,32'hc7c10005,32'h8fdf0006,32'h23defff9,32'h0c0001ff,32'h23de0007,32'hafdf0006,32'he7c10005,32'h46001003,32'h46030000,32'hc4230000,32'h34210030,32'h3c010000,32'h46020081,32'hc4220000,32'h34210030,32'h3c010000,32'hc4210000,32'h3421001d,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c0001ff,32'h23de0006,32'hafdf0005,32'he7c10004,32'h46001003,32'hc4220000,32'h34210030,32'h3c010000,32'hc4210000,32'h3421001c,32'h3c010000,32'h45000011,32'h4600083e,32'hc4210000,32'h3421001e,32'h3c010000,32'h4500002b,32'h4600083e,32'hc4210000,32'h3421001f,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10002,32'h46000800,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0001ff,32'h23de0005,32'hafdf0004,32'he7c20003,32'he7c10002,32'h46001803,32'h46040000,32'hc4240000,32'h34210030,32'h3c010000,32'h460300c1,32'hc4230000,32'h34210030,32'h3c010000,32'hc4220000,32'h3421001d,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10000,32'h46000801,32'hc7c10001,32'h8fdf0002,32'h23defffd,32'h0c0001ff,32'h23de0003,32'hafdf0002,32'he7c20001,32'he7c10000,32'h46001803,32'hc4230000,32'h34210030,32'h3c010000,32'hc4220000,32'h3421001c,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h45000017,32'h4600083e,32'hc4210000,32'h3421001f,32'h3c010000,32'h46000801,32'hc4210000,32'h34210032,32'h3c010000,32'h4500003b,32'h4601003e,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46010002,32'h46011041,32'h46030842,32'h460418c1,32'h46040902,32'h46052101,32'h46050942,32'h46062941,32'h46060982,32'h46073181,32'h460709c2,32'h460839c1,32'h46014202,32'hc4280000,32'h34210020,32'h3c010000,32'hc4270000,32'h34210021,32'h3c010000,32'hc4260000,32'h34210022,32'h3c010000,32'hc4250000,32'h34210023,32'h3c010000,32'hc4240000,32'h34210024,32'h3c010000,32'hc4230000,32'h34210025,32'h3c010000,32'hc4220000,32'h34210030,32'h3c010000,32'h46000042,32'h03e00008,32'h46000801,32'hc7c10004,32'h8fdf0005,32'h23defffa,32'h0c00016d,32'h23de0006,32'hafdf0005,32'he7c10004,32'h46001001,32'hc4220000,32'h34210032,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h0800016d,32'h46010001,32'hc4210000,32'h3421002a,32'h3c010000,32'h080000d1,32'h080000bd,32'h46000801,32'hc4210000,32'h34210028,32'h3c010000,32'h45000006,32'h4600083e,32'hc4210000,32'h34210027,32'h3c010000,32'h080000bd,32'h46010001,32'hc4210000,32'h34210028,32'h3c010000,32'h080000d1,32'h46000801,32'hc4210000,32'h34210029,32'h3c010000,32'h45000006,32'h4600083e,32'hc4210000,32'h34210026,32'h3c010000,32'h45000010,32'h4600083e,32'hc4210000,32'h34210028,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0000d1,32'h23de0005,32'hafdf0004,32'he7c10003,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10002,32'h8fdf0003,32'h23defffc,32'h0c0000bd,32'h23de0004,32'hafdf0003,32'he7c10002,32'h46001001,32'hc4220000,32'h34210028,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h45000011,32'h4600083e,32'hc4210000,32'h34210027,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10001,32'h8fdf0002,32'h23defffd,32'h0c0000bd,32'h23de0003,32'hafdf0002,32'he7c10001,32'h46020001,32'hc4220000,32'h34210028,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10000,32'h8fdf0001,32'h23defffe,32'h0c0000d1,32'h23de0002,32'hafdf0001,32'he7c10000,32'h46001001,32'hc4220000,32'h34210029,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h45000011,32'h4600083e,32'hc4210000,32'h34210026,32'h3c010000,32'h45000026,32'h4600083e,32'hc4210000,32'h34210028,32'h3c010000,32'h46010001,32'hc4210000,32'h34210029,32'h3c010000,32'h45000050,32'h4600083e,32'hc4210000,32'h34210029,32'h3c010000,32'h45000074,32'h4601003e,32'hc4210000,32'h3421002a,32'h3c010000,32'h4500007e,32'h4600083e,32'hc4210000,32'h34210032,32'h3c010000,32'h080000e6,32'h46000801,32'hc4210000,32'h34210032,32'h3c010000,32'h080000e6,32'h46010001,32'hc4210000,32'h3421002a,32'h3c010000,32'h080000bd,32'h080000d1,32'h46000801,32'hc4210000,32'h34210028,32'h3c010000,32'h45000006,32'h4600083e,32'hc4210000,32'h34210027,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10003,32'h8fdf0004,32'h23defffb,32'h0c0000d1,32'h23de0005,32'hafdf0004,32'he7c10003,32'h46020001,32'hc4220000,32'h34210028,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10002,32'h8fdf0003,32'h23defffc,32'h0c0000bd,32'h23de0004,32'hafdf0003,32'he7c10002,32'h46001001,32'hc4220000,32'h34210029,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h45000011,32'h4600083e,32'hc4210000,32'h34210026,32'h3c010000,32'h45000026,32'h4600083e,32'hc4210000,32'h34210028,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10001,32'h8fdf0002,32'h23defffd,32'h0c0000d1,32'h23de0003,32'hafdf0002,32'he7c10001,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46000801,32'hc7c10000,32'h8fdf0001,32'h23defffe,32'h0c0000bd,32'h23de0002,32'hafdf0001,32'he7c10000,32'h46001001,32'hc4220000,32'h34210028,32'h3c010000,32'hc4210000,32'h34210032,32'h3c010000,32'h45000011,32'h4600083e,32'hc4210000,32'h34210027,32'h3c010000,32'h080000d1,32'h46010001,32'hc4210000,32'h34210028,32'h3c010000,32'h080000bd,32'h46000801,32'hc4210000,32'h34210029,32'h3c010000,32'h45000006,32'h4600083e,32'hc4210000,32'h34210026,32'h3c010000,32'h45000010,32'h4600083e,32'hc4210000,32'h34210028,32'h3c010000,32'h46010001,32'hc4210000,32'h34210029,32'h3c010000,32'h4500003a,32'h4600083e,32'hc4210000,32'h34210029,32'h3c010000,32'h45000074,32'h4601003e,32'hc4210000,32'h3421002a,32'h3c010000,32'h4500007e,32'h4600083e,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h46010002,32'h46011041,32'h46030842,32'h460418c1,32'h46040902,32'h46052101,32'h46050942,32'hc4250000,32'h3421002b,32'h3c010000,32'hc4240000,32'h3421002c,32'h3c010000,32'hc4230000,32'h3421002d,32'h3c010000,32'hc4220000,32'h34210030,32'h3c010000,32'h46000042,32'h03e00008,32'h46000801,32'h46020002,32'h46031081,32'h460300c2,32'h460418c1,32'h46040102,32'hc4240000,32'h3421002e,32'h3c010000,32'hc4230000,32'h3421002f,32'h3c010000,32'hc4220000,32'h34210031,32'h3c010000,32'hc4210000,32'h34210030,32'h3c010000,32'h46000002,32'h03e00008,32'h46000002,32'h03e00008,32'h46010002,32'hc4210000,32'h34210031,32'h3c010000,32'h03e00008,32'h20010000,32'h03e00008,32'h20010001,32'h45000003,32'h46010032,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h20010001,32'h03e00008,32'h20010000,32'h45000003,32'h4600083e,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h20010001,32'h03e00008,32'h20010000,32'h45000003,32'h4601003e,32'hc4210000,32'h34210032,32'h3c010000,32'h03e00008,32'h20010001,32'h03e00008,32'h20010000,32'h45000003,32'h4600083e,32'h08000000,32'h68010000,32'h20010000,32'h8fdf0001,32'h23defffe,32'h03400009,32'h23de0002,32'h8f7a0000,32'hafdf0001,32'h20020080,32'h20010080,32'haf650001,32'haf620002,32'haf610003,32'haf630000,32'h346323f0,32'h3c030000,32'h23bd0004,32'h23bb0000,32'hac250001,32'hac230002,32'hac240000,32'h34841f86,32'h3c040000,32'h23bd0003,32'h23a10000,32'hac610001,32'hac640002,32'hac660000,32'h34c61f2f,32'h3c060000,32'h23bd0003,32'h23a30000,32'haca30001,32'haca60000,32'h34c61f02,32'h3c060000,32'h23bd0002,32'h23a50000,32'hac650001,32'hac660002,32'hac670000,32'h34e71e60,32'h3c070000,32'h23bd0003,32'h23a30000,32'haca30001,32'haca70000,32'h34e71df7,32'h3c070000,32'h23bd0002,32'h23a50000,32'hac810001,32'hac850000,32'h34a51d32,32'h3c050000,32'h23bd0002,32'h23a40000,32'hac240001,32'hac250000,32'h34a51c8e,32'h3c050000,32'h23bd0002,32'h23a10000,32'hac810001,32'hac850000,32'h34a51bbb,32'h3c050000,32'h23bd0002,32'h23a40000,32'hac230001,32'hac240000,32'h34841b62,32'h3c040000,32'h23bd0002,32'h23a10000,32'hac610001,32'hac640000,32'h34841b50,32'h3c040000,32'h23bd0002,32'h23a30000,32'hac230001,32'hac240000,32'h34841b03,32'h3c040000,32'h23bd0002,32'h23a10000,32'hac640001,32'hac610002,32'hac650000,32'h34a51a94,32'h3c050000,32'h23bd0003,32'h23a30000,32'hacc30001,32'hacc10002,32'hacc50003,32'hacc70000,32'h34e718e2,32'h3c070000,32'h23bd0004,32'h23a60000,32'haca40001,32'haca10002,32'haca60000,32'h34c6185f,32'h3c060000,32'h23bd0003,32'h23a50000,32'hac810001,32'hac850000,32'h34a514d9,32'h3c050000,32'h23bd0002,32'h23a40000,32'hac610001,32'hac640000,32'h348413b5,32'h3c040000,32'h23bd0002,32'h23a30000,32'hac410001,32'hac430000,32'h34630846,32'h3c030000,32'h23bd0002,32'h23a20000,32'h8fdf0001,32'h23defffe,32'h0c002461,32'h23de0002,32'hafdf0001,32'h8fc10000,32'h20220000,32'h8fdf0001,32'h23defffe,32'h0c002461,32'h23de0002,32'hafdf0001,32'h20610000,32'h20220000,32'hafc20000,32'h8c210000,32'h20210000,32'h20030001,32'h20020001,32'h3421008f,32'h3c010000 };
endmodule
